��/  ��^k*��A��D@7�քW�g̝�G�^�T�|�IVϪ�y�p;�5��p:#�oj#�_��J��≶���j������f����v��X��#Ο1�v�S[�T*]ZZ�'��b�&���\�uQ8)����/3{���>Bm0��̳>���T�d��#/��[r�I��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P�A���1~�-CtP����2۪AФV�_�L*c�ƿ��z��*6u��`6i2����>T�$� ��M}���rSf�8+[ϡg*�B��ʲY���?GL��-ʥb���$ePF���:Y��U�S�ؠ��!�~_CXmqY�����x����E�[<�*>F�����_�דYn�C]2I�E����a����]K�?6+�?����)���j����F]2uo�Ŏ��\���S���GP/y��A��gr�� n"/�� ,���&�x�M�����|f#��v(����(��ٴw'֟a�m
��pۋ���U��I��}��ZT�l�:7��\��?ԗH!G�}"�$�ܖ�q[�hwZ�
����[���*m~Mk�{�H�
>�3��f�9,sJF��#[�pꔵ�b)��B+��k}�#��_�C
툍Ъ;;�At�(�BU��, u���R� 7��-�]e���+_AP�u���L��|�, �A6���D�wP]�?�m����naҿ�[~B>m��)���&�-�Be����vث��q�9�#��L��!���%P6Ҫ�/�d��c��+
~���
w�ϥg��f�{�A�`��.:0�wG����lR��l+���((\V�U�`]p�|"X������9ٱ5�M��'.W$�'�i&��QoV�rj��"'�Lq5b��[�WIq �J礣~xߎ��5e��?*� ��j�;�k�=��V�o����D6��W���ֱPϧ	��wa_��j}t�|��hꯘ�t���
@Z�.�*?���2-��u�B��:����0�I3��A��'�#�]Ҹ����9Xdx�$È|�����/�w,I=�g�G��CXE����k~!L8��j1��b}�4_wOY�-/qj�*y*/\��DX D�9�� �l�-�	*��Ķ�}��g�!�D̮�0��TX�^O:��;� ĚgG�Lg�o=��h�C�3�����;L�r��N�Y�B]��;Ū��0��������8%��h�17��a(4� T*38��n%����e�͏��>0;(+D�$�V+���j�}��(��
��SȐ���[��b1�J�)h��2p>�V�#08K�;�,��a���~�zT�xz�[��>L�3i�|=�Ҧ�*V4��m=4��[��V`I�9�.r�E4�%�d�B��WM���d+��V)��<���ч�����G=���^o'7����[Q���䰪xT���w�"�����a����t�$�����	��2�j#�/,��E's+jx	�qӾ1c9�/e�C������R�=)�{����D,{�:+N5�TI8zK6��r/ �kJ����jt�M@#{�ߓ� ��9_��`d��g��1��5d��c�f���	�� ��
���e���.�D��">��w�U��%[;�7��������������.TL��;Xǅ/3g�+R��fL/����+��O���j���;��Z�����8(���~��N�3.@�F�iH@�]�v��RI��ihc^��\{�ck̐d����P6�{�!����	B��7�1��@)'ō�߸�-�1��kǈ�a�v/3���$�P?O�����W��e�X���H�y����aS�d�� 	i�ڪPR��5΃�
��N��{'�4�����%}ۢ���{�V{�s�41��XX��e1P�lu�ht��:o��k�OZv�S+��4�%�(��7��a
����ʃVG�N��[���*ė��Ɓ�ŕ_�T�y�x,[�uM���9�����7BjK@��G�� �f��^��b����}b-���.X�߽k�mrŭ���o]������ܤ)C�)��P�N��gQ�n���?���*V���"���pc{r�����õ/d�^��s*�Za�a�I�T�b,T/*�d�m���(�Eb��J4�ﲗW�Pvt����0�c/_���hMʿ��C(^}w*A�����F�<>�	+�a�j�S���H��N��pɭ�0�FC���n�F�>��ˮ��Nnf�@I�����jzL�dȏ�Rl��Q	jF3z��	�W��u.iQ�O��.���; 55����cwL�0Y�NDj�@�z�HI"�~&�bk*!��a�P��=]��^͡l:�_~O�o�UG�)���^��UI<��+��[�� �<���I �/k��,� �s��'̕d�� 3t��;z��Al���aO��L65�
O�M �|����Ǉ���1��k'p@����%�����*�O���x��Ϫ��S�,v��fSX2��ªΎ���S/��qK�t'��~��+�F��v>��\l�R::g��2=pM��>��Ez�<_!��U7W�Ecu<aM�|��V���3T\V��ʞ��!y�5�%�X"�\��&�W\�7i��ch����F�̯[yG�t�����g�c�sp���׶���L|���S�c��/���ǙS�13D�ͻ��p�Ǌ/#&l����WS�b�5�IٯN��A%�b��ӌB̆Us��D�ʉ^E1��[�%M]2�J5M�%�/J�XSO��ڍ;
z���4�D7x��J2ʧ�i)i�)��>�Ȑ�[��[u��/%��By�����-�a{�a`HKL�9
SrUYd��%�k#ߟ�dr�S�n։���3���*��M#h?
�,�c�����/��7Bi���K��<�U���i�A�sMx�FisŸ6�!!�AGȂ�a�I��c����J���t�tg��n��Y�S�i)��C��؍��� 1��6=eڒ�p��05�y����x4�|���4��9k�tu����]�^Jmz�d
��6,Kձ��h2�΍K!qO�dߚF�����e!�.��)`�b/���_����oΔ��\�� ԅ��3|غ7�G�=� ������>v3��ڈ�폆�.�{?i�z��z��IWE��G.M����۠@�oY�2��	DAa��'�h���'-�Rێ�		Q��S��$��/����{�Q�v�	��D��T}.O������ ���M���L�#?VHs����dx�D?���8�{WcȐ�2<�$4e�F �/��N}E����H�| +E�$
��.ݷn�WH�
0�y���:��H(�@�������]�-�G0�~����<�9�سb��T�C�(��~���<~��s��\2VT54�����&�,ju����a���	`��i��K�2�.[��QO;�f;5�X��vL7��3�z܃��r)��ٛ-_�w:�\0�o�f�/�JS��V�Ce��GBi��-����ym�����I<���7u�ϥc�y�ߦƪc�}�n�j��/7L���7��J	��w2TX��pT^�X�o�H���r�k?�� �t���x:��~���X��gB����;�;�>��2��S���\5m�)��fE��JP�����HP�rb��
|��?���Áz?�4cD^�~
�Jl�9���[`����c�� ;�c6������D���K�FH|�tۡ�x���[�w{G��9���]��r4-��a���
6����㡙\�
P�s���5v�8�;��������r{\����+�;��[��kT$e�C�B"�މ.ȩ"(7�P�^���3�F�L�3�gv�������Q�wf%�T*#S2GV��FDِ���1�!�RKg�����+��\��$��'����t�����y_r��,�;C�����Oqs�#)q�j~�e�~�F5�|'s�m
���?�����_����������>�� �i���	���TP!b��=�<��z�k]%�:��$��0��-����sq�=��7����|s[���`;�_�#������ϴ��5�<!):j�G��a����'����M%~����?�9�<����|�@�b�Thg`�y�����	< 2��8��5�z�:�K�a`�~��xH��?ag�Y3E��M��n���n�eC漲20"�bh�gd!�GQ���Q�,��ע�yz� *�ks���S��E�E9��X`�d=䡲�Q��W5j���c�[ۀB��A�6Q������Ek0L�6 �Q�z�mB0ݣ@�D&W�Nt���l@��+�b��ѵE��է~���T���U� I4�Qw��薌�.���3׾9����5u�n�������"5������q�������I�Y�1q�����%~x���ĽJ��7|%���kj�$sL���m�(���qܣY{S���ul#�q֟��� ��%��/�	�M
���UT/��# �O4/v�X�'�.͍�Q^�!c�4O_N	7�M�<M���mrm<����a`��+{I������^��Q��U{)���B�Ƞ;�i�F�AaA�(/s�EjL"�1���J�m+�n �!)d(�����u5�t�����\?��ռO#\«��\����3Uqzy4�羾��=�OJ3��f��ʫ�+�����̨r�\��`^�S�D�^b��Ꟊli%�x�I�P���1�Le44Tt�~��`�B=~��b;azs�=č��#�/��U�g.l��<�I_~�Z��p@�P�*L6�u��[���@����|{>\,-r�46��R��v��p�_|�A��f�PȌZ�8�&+�BYz�T>�(c�dC/�0Tm��K��2Hƍ� �1}�����6)'<�OY����R\��c;���;�t 5��{i�g�����e��*:�{���� ».�:�� ,[��%�%?����̄a�bS7e����.
eeQ���?�[�Q��Q�c|&��@���I
��#�X���׊m/�-�3
֖KO&��`OG��H�_����s �c@?5���U"�J�օu���"N��6�}��:��"}�X��Hn���5d[A�?��
��-����n�
���<�N���B�ȑ(
�����`y?NU�6�V4�S���� �17L.1�}ϥ�ß�{�a�^-GU�A ��u����o�~؜^��ڲ���J!�����|D-�ҽgms���+��4L7�C�S�V�	�#!sxb�Ҵ�_ڄ|��"�ဨ/��N��]�ʅQ(�Q|��u߇r�p�?f��=ͭ�Q�%�G�Ȧ��:�V�xBԢ+=��o�o��q{�'}xE�)����)�|aXD��>����k���GLDɵ�7��)����ȸr<�Qk��q{4?�#���r�m������V�����	����^?�xJH�y�Ϩ��Sn�/�<�$�Y�R�\r9pG�܍�� ̵�WLs�4B�:�#S6Ĕ*V	���2��n�c5|Q�>���m�ԞL�ܡ�ƕ���>z���l��h���f�@�����5v�M9��_�TF<�u3�u�1:}�W���M�T� �ٲ�}��9�����}c�/��yNms�I����L��}\%p
�r��x�~�ǋ*��K����@�d�_�]k)��ܑWO>¥BT�I�=;"Ǯ���|ǟ��o��	� <�\�$4��*�(7��%��C%X��Bw�Ә10����|�����%�J�{��^}�9ׅH�r%7�`�Ķt��z_�9�'	��2m��0�?��=)�{�CN��t@(�����<۲X1�4�%���r�w���,�Pⶮcy�푎FN��<��,A��y
BI����]�jdY�$q5.�˖ڧ&���WmI��U�b������\���u=�RHtv^�ي�m�+���6������S��U	z�J�nJx<�t����4g���(��>��}��d�&�~e�[o�@��MU���:�]Ȣ��/T��L`b#y����)�֠Gu�U76��Hr(�]��8��)���sN�h<Xw+�q�C����~�Y���0�3c�8�R�T�1�\��c���k��S�L�}��%�a���ڤP�K������h�+���V_1���6��R�)\��}���f�X�t�,��m�g[S
nv����@����E���/[ ��N��GbL������:�Ti	�W:t��S������u,���C �w q�� D+��
T�)�y3� ��!p���IFRs�.���\�H����L�Q.�=�!hS[I]	
KL�R%��<U����*Yo�
�(U����To�@ei�s J�

�'�6�����M�r���/Z=���z�[ڹ��m�����[��!֭��( B�^'�b&�����:�� yKB�h���x��*���zJ����ĺ���k�7(��̲����Ms�/�s�b``N^�)�b�G�3<���|����V�~��ϝ��hFB���|��h�,%��|.EU��>���%�}�}�u�`��M�xɊ�@a�vvj`�e�g:��x��j�n�<�.���(h��<�J�7����� {�9��3�@��zG0��ٛ�Bul/]1�;|6*:j�r�(��I�+�<����!>F��mD���2⣀T(>�O@��������<���cQ��\߆"3JV��b<Uc:��:�#��{�� ~�of�~�,�ÿ?�w�FI�(d����ShP<1 ��`w�f���&���b��:n+��y��W�1�}��f�_����[#�=���>x�e}�bs�{$ӸŶh�L,�Q��U����9_�^���3��~v�}&�9�/��?|B�:XY� x�A��A�?�j�Oo�+0�+�/��;���}=N;z`�CKP�ݾ:�H�Y#���	��q��͸c���D,p �Z��#4���o+�uk�,��5�� y�����`Iv&� ���/nC��O�f�x�ʡp���#�ݦ��Z��f4���ƫ�T_���@�'�!�ca�	�}���v�m羪�(]�Y�fM������-�=s�)�K��6.��ͽ�#���C�����#���ri��I�uL���(�R�q����m�u-����3!<#�@��@�����!𰰝��m��A��0*:��Z��K(�&K���L(���8&Ix͂}�/���hj>"����<BW@^��V>=��ad���?�$��J�$���~/�:����+��S�k��������fP#��#�"9�$���am�!3?�fBJ�&E� �$X?7/Q�|Gy���*����{t�N&��Jd��f�����ۥBD�9�@��]��~�y$�0��v0�y��f{��[�=&��~��K�x�~y��"%!9�ɱ�\ha}Vu�/s�N�~���\��R�]���Ŧ]���ؘ �Yt�J���%�?ױj�1�6�J�Zk[��i=�9��7��U��E��l'���33�t�(�P��d�mQif�y �
ǈ�~�J���}��awcuhQZ�m98����Y����}��Zؼ�Lb>T��o>q��f�{�<Bf���k>�[���������j�遆�ۼ�U�.��G�"��O��q{x��\��c�m���꽥�LqE�X�d��Y�Yq`�f~�� �O���7�:���7�ۉ�-gIex�[�_��{{	6"[i*�[�b�r��)5@+���Wv}�v�z�V��W�T�5G=@�;����>�D5�V�"�, ��*;��4-��[ޑ�h��`���*uի���lv���e��-�W5ʼz�<�W��o�P*]i$��f��Z�S��V)��dn��}gE1J|Ҽ�.��'0�_|�����N����٤m�E"�@J����Sv,P"���5Y̛Dዙ)�.�=�� @"��m�4���c��)�L�ڟ�q���B@�x���ܕ]��q�+��d���)l75�3�U�q����?��n'O�u�U�L����8�3�(e�ɇ҄H��LT�6��[�1o�z���ub+U/S�Og/uX�]�U���Ϟ���]֭�x-�v��.B_�+^��XE@�̿�gL�"�j� �OZGk&���Z�[�l���Ч�q���&bksn���Zy�/5wI����^+��&0X���I`
!`'S�TC
��X����ne`��u�~;�ĩ�W<;�D(�����m���t/m-^������7J�6q'2�ی�����}�lg(�.��Q�����n7g���J�̍��U-���J'�%&Y��7Q#��*�]��EM�V��K��IW��DX����y�,��]���&�D�ٳ>dO6����K}�˻-6PԲ|��s�1�x���s��v]M��VףjjA�K��q���!{���|�ߖ5�)���'�7��������(*n�>�A��Q����5{XN�7��e��af�L�e����}����hNʜ���Jv�t��f��D���jiF�w���ȑT
� ���>Ɩa ־��MN���_���q&w��7�15�� �D���#�����8�ҋ����&����R�?����x���������G�]�2�RK#�g���~"�~Js�,�Yӕ]*�@� ���	kE����Z�����\���|�h�Ɍ�Td�i�*��g�
�wYz�;_��sq/m�.��v{;t�seM�7��l�B�eNھl���W��B�X.2�y�1R���~�7�w���OՁ{Mu��)��)?�%+Y�B�k��TsAg��6U��ָ�wA��S�f1�t�p���_���;b���J-?���T_������M��`����SE��6�Ä����;��D�$_5���#_Ul:�d��<`y��6��g�U8���]J��c!�qL{�&���qz��Y���׺b�p�	����O��K�� k}y'��K�4�_'�����i�#��$�7e@��x��wg�,�|��YZ@��Z��^VS�XSS�Ps���H���Q��8��m�j4o ����v�t����;��՛�,\O��:��]?-U	��9_3(��Gkaf��B +�ߊr4����C	������
�E��i$C���CŅ�&@� ��'k�Bz>te�-%�����KH�_j4�3��Vq�'ͥ@8��\��3ѱ䔒����n�KDX�T�[e�qW���ݻG{�OѺњ��!�#��4�{��f��G>�,���r݆������2�u9�\�#;�9��Y����ol�r7bc$�'K!<e|̛Y�i���dV��*a<��?�/7�	��^���4�ĵF�1�SmT�����P�8a��sP�&z~��H2��7��-i㶝���B�&�m��;����I���M��T:Y�46��$�oN��7yȖ�qn�U���=b�}J�Яe�
iT�Ў���n�G|̞l��"H�F��'�c�]*�L�dA�ƭ-E����|)J��S��.�~^Nډr���{$���"	<�T��K�alQ�O�Ԛ���N-�j��D��1�5�޷8y'�"�|w����=b��BS�]!��v~�=����m�J�+,u�V�9�؋�?D�j"g헺�}���xW0�`٘��:�G=�$�J�[F�������7�������i�)p��\�L�bf�qy��#w���f6�f;T8�������)~�pТ��	C�C����q�(�������&t<��!�	�Z1َ��PY�X����������u�*�
�]�ĦX��n��Z�̶y��G�.
���n7k�qB��y�W�:N8ԕ���oۏ�>u\�Z���?{s`��9%��I��HAJ�ot��0Vּ֊W��.�ە'X���6Ju�;��ri���:��ot]_�MK��^����b�X��iܺ������Դ�I�Ԣ�>�z�H�f8f�9��yZ� �5Qs���q�R��xJP�K@I�5_(E�*�AUw�Q�1&�D�
i���Nsx��hevyUX8ʐ��_!N���YX�zs�&BRV_�k��a|vA�E�7���4y�����7�#�o�.���g�����+�S|S⥣���a-�1rt��#-�R�XE��x�0Q����E���=�fS�9E�[��߆��Y-�
�oB�3�ɴޠ2��K/G/2$K��5<Ob;���XH����w:z���(|��0.2D�,WRmz���.�Jz��6��~@���,FUfdƹ�_�`��W�W�Z��-$��&z*#è�4��&~����u�M��d����V�v�dj3g���Ȏ��Z�=��I����yjt�pf��=:3>�\G=l9���Th� 
�*��p�"��B��:�*����l��L�ѫ��i ��U�%Y��tv�""i���bA���~�.�*�ؖ��H�1h�ݷE�|�����=h��f��w�=vb�U��|K�W�ŷ?�*M1V'{���
��Ń��F�j�A�*�[l�#z]p$#��so���p����+��J��;�K�X�S���1-���j�CPhN�*N����o��ǜ����<Y5N컸�⌨  U}2Pǡ�aX��ɑbDE�+\��M�2�̓s�a�цg��	��Tl[�'Ks��&$~���e�be�B�s}���h�� � D����m��fM�f�U�|��vXc�
����C5�ν�p�P�©Ɣ�UU[PM���DO�X��k��q�Y�7�qi��׺���&����,�ws�}6�V^�g%l���`)�R�>�^�����X6W�-=�.J�iX��+c�\�!/n��:^ay�B��65����u%T1���i �Y&� ��~��Xஸ	�����O�����`�z���=�9]�`����PR_�5��L,e=��b�&-�&f �dY�Y��8Idt\��s��9��zhK�,9]�IK8�����(�|E|r�j�`�u�חݝ�.F*PS�x���f�ҩ���pf��a~��J��k��M"&�}Q��l a�`=�'�9����+jс}��9)�LT������U�̢Z��+N^��෎ ̀�Ŋ׺�ﵺI[P��~*��PEϦU��pB������z��7eŅ����U����$ȁv����y�����n�l|N��Ʒ��a�-��W��S��Ύ+���$$��R�9jo��"=iʺ�R~aWK�m�ndz�)�s6��#^��P�;�E�:�Ps��_��y��ð��1��a�_ڈL���z���F ����r��7������a�g�
�����p�[HMz\"8��p�
��XxH,UGCR��Lo�+h���=��Fa���ɺ�2{h������5�q��#��}�V��;;���5�_&����F �Z�D�A�ӗ z�C��|�ë�W/���[�|z.Jь��A[ٻ��*�'M0v��D�ko����g�F)0̈́_�_������݈M�x�?uC��C�Տ0��zLV�у2�9�}�ɐћ�:�w�i�>�+.Y�vݘ�:F�̰�ܒ��7�֓��,�eAAc�wd�C��������V����t�w�uF�Q�ʴ�"f�zzY��I>�����:�6��L�_��!�,�Q�y����e-��X��xPf�0H�X�*[Rˑ��ރ�Tk���DA��'������3�E=U�R���2}My��LKȔ�0�hd�vE@�k�|����v&����W�w�#NI
bu6t��Ef0i��(VV�L|]2Y�3DST�H���$r2�V��M!�x�L,��cԚ6>P�n<2:��l�'��%`Z,���;g*��$ �:��R�^�����E��)��7��!�-������9�WΠƧ6�CS):��;6��"˓$�Ux�eX���k	85��񒉈?h�-`��@���Gd}	-ݸ�g~��"	w�E6�
1ErfJE%`5q"z�<���?�׏>�$
V�nZ��I����I NY��X+���h�׻#S���F�iv��9�;����|U�&�5C��]��9�7=�h�.	Z �p`��)Q�u�J�+6$�)�j�CQ7γu�s��J���V�k-����K.s|��1��~��(���A"�4�@[lS��t����ț�n#!}�U��S�&��O�D���]�H��_0�1��������4+K����]Fñ"����<HY8u��<��e/����o�i _���G$��q�v�'z0�4*�%o21��̂{t�,*����p��}9���l�q�0f��]��/�L"�jx:���0"=���g#]d�d��M���3�8;�DJ'Hg�f]O-��W|��s[>�w�Ms^f��<��[�`:���c!r��U�7I��+����1�`O��IV$�@5_*���������+K����?���:�>��hؤOU�:4�C;�r���O$� ��-7*=�9Dd���9{�@U�Ƞ������8.9���e�A���M� �%��<��;3網��(�l���v�m�X�wf�Pj}�����!��)������˖k���)�H�K�C2�}�/'�o�<�l����⽋��goO~[�3�ե=� w��%��N%k<�Z{��7%�.��X5���@^�[��2/�/����If��y���ze��xG�n�prF�����{>5��	Rˍ1�u6�hs���۸qL�:o�%!J��`&�ʈPg~TQ�ـ��W�`���Q��&��2�����w<����:�JYgO�Фb�0��0���O�],&ڭ�����o\O;3�.���эU�-����M�4���YD�7��R%�j���BMsƱ���,ۻ:�AD�a��4{��3"�����!t�	�Zј���g;ކ򊹥9wf���3j���j]�5<E3s
�Y�W-�Ϯh{/��}V-F��f�y�wKB�!4�[���stC�%�A���8���(�О���xR�^:��C�V"�Ap���p�Y��8S=O��W(Q6�4P�;M(	����Tx���(=k���^daV�9q:F]o��zg�s�+�$��e��mθ�������O�����}�%�_����шYKc-S&&�jאe;5S�O#4R�u!ûd6���a�G �Ic����eD����HJA�`N��!DA���X�>��:��d"��s��Àh:�d�����2j���(�@����F��H~%��A��9��(�t��Lz�_/o� (8��%	��3���͵R��R�W�Q��M��9T�M�-b44�ɥW�gA1��ȿLS�#$��Om�nV&�wV#�s�S�D�8Lݜ�w��>p����%z�=�=�A3�G��Kx��O!U��8�Iz�<5�S���7 _�gEgw�=�IuB��S��W[����p)�YӼ��{��Ji#Ќ���x���)URFT�-�e�x&+;D9�5IF��9CK�t5��
�6~	3��a���E�s��rujtj�ĞlT�0�b��m���E�4�Ϸ��dU�8�5`PvC��#2���g�EtPI7�Zm޹��v�m�ki��@���D{��˳����@?�O���zm��r��`�wT�A$����ħ�~f�P��`<5��9G�����I �9}�o~]#i5w�'�� Sc������&��lҧV����\�17M9�[�Z~�����������//�o�i��Z���t��a���i@���w����&?0~�bgn�#�F$���B���;䂛ۋ5-��`N�����٘;{���=NpH��Z]�_�K���=v�b��aز^&Hؤ��y����W����B�8�;#�k+��㢜?XN�f� �k�Ȁ����GGGd3*��>�~�p��S�*���2��=F�H��8GH}ݴ�&2>���׫��)Ҝdw0��幄@<�CD�P!@�p{���GSH���%Q��h�b�BR$/�g���\:u� �@S�kU��PQ2Z�b�D�B�z3U�����0�R�]��z>�QR�Q|����������c��Cl�[3
D�7O�Vdͯ���~�/E}�4�Ayrǎ��y�k���e}5�#R�=�lH,(TF�/S�|$������Jȼ����F�:f���/l5�0�]a����*��P&{����m����Q�.�����Q��j��O�+��	�oJ��wX�Z��@�v��E��K�*��U�����:�����΢����=��^����Bd`�E2?��+
5�� 7`�"͡
P�ފT$���� �_���B�H`r�i��fAȰ5rn:
;����SB���K�2�3�_��F+|g��~�,��)��Uj����&��d.b�9U��㢸�	kzR�_)";2u����8�WYDBk�-0��YZ?��� 
�����mXǫH�!�>ݤڪ+��y�hxt���.w��7i!#d�8�̑g�)�at7���d�^?�^c�f]�_�8�B��(m��93��rt�C����x�jl(��0� 520��B��r�й�L�f��Z�=%�?���W!�eE�jY+ !���]G�y����Ǯ��J�v���N���>+��K�IBο����8f���$p�3D7�����O�� F^��X�ѱZ��Z8�F��q�x��% 0nx���)i�Oht��A(_bza�,3EQ��]!;H�d�-�+҅�BXvcx4�f�&:�����s�H9��0�E8
�����NU�X�+���2��h���y�y�O��(�I����Xx��9C�C�l�f���e_�������Z�N�%�e-R�ً��;�v�;o_���,�2��5.�蠬B��4R�o�
�U�2��T���b�]���� {��ۃ��ė���f+O��pL�����2X�`��!�޴
��=��P[j�k���$����L����בm��T�>�զ�f�l����M[�{�]]�	iá�`�A+�Glv٬���1*��j��R|z���n̃��`��o�V���v�}KկX�/����BoەqG4Yu)�.p?ˠ`�'���F�/I��v���(A�L��$�w߮Χ�;����LȀ���ׯ����l�Q3�DD�,	�s�M?N-�s�
(�ZNҤMI�w����32��Y(2D�z�ɥޗq��&]��M�1oS�
�5"��&��xM`j�xI͖��X�0_��2:���HA��ԋ���[��*� �/�5��1�d8�)��	�o�/tfYe�pX�ŀ�uݗ(w�0@_�^6�����OS&���`n���R�@�8��k'�K!<�?�F�O�A�`XKo�B](g}��n� �5�^���b���Oe�"�]D����\��/�r�QL�
-��T��wf������[҉-�wxP��o�7k�#ơx���Y�ա�3y0T�v}ߍ��G/��k��Q�3��mqu5!D��L�5��`(uЁx>�*���~�3�E-�y&*~�gm�߆&P�K�h7�VL-��/�^Y��{ E'�9�&��ho�Z{	�Ԉ *��X�/�J1�t4k�2�͙�W�-����� �}����%��� -�@�d���,��.p2�*׳��ȿW��%.�h�U�(����M�2>0�r�z�O-�M���4���M�k����nB{��h�	��7���)(XG�Ww��i���S??���$�HG,G��=6�bz��X��z��9X�5�p�S��͙��W�E�mo/|�����pH��4w�=z'F���N��_l�~v�=�GOE?�Kh�ct��qМ�ag'� 6O�i�����q&�=�/��i�� �T�0�}-2v�"��zk�f\}Mbo8HP�Im�t�ZzL:�����:`�Lbi-����������ZDA��|g	�֡��*���:-Y��Y�������Os�T��I�!�^�:&R`���C������M0�3t�T��)���&ߞo'��@dظA��Jyƥbɀ��Ol(��4 �yqm�2["� H!E�}s�l�VXD7�����"��JE!a�b%�9���r��W���Yx��� Jr�bIMA����x;����<(�v'�hѵ˓��M�W� �)8����-?]S�Y%�9�+��Չ;5�J%��? |#}�<n����/0,ֺ��30P��NY��ǲ�H�v�{@��h�N3[َ&%�bf7Z����$4��ا����i��I5�����}���T�0z�����L(��������#'~��J;������mh�������m �`��7s����t-`=����!�n���\���f�FK:&���
!`����嚺����������b2����끙UgTSL�rRC���9�=(����pk˓����8
)��eULY$�;+<�B'\Dyq˦�+|��u�x�6@����"#���B.i@kJn�KC7;���]��X?(��uϗMqM��!�T����gQ³U���Z놡�Z�^h�m�}D��`�/�sEO�E�XŬ��=2�-���Z]��5]�=�n-�Y���Xsc�TH�����a)h3UGci:�����fa��eg�eI�u5�n���p��c���.�t.��1��5|�7"�7A�������/�g�C$��{'��d������l�-�w?�m��}�b���_g[�"2v�%����ۚa�/`<�����B�)�Ʉ�s#�mモ[��݄�s��Kq�0q�ٻBo�P�R��Y��Q�8����j$#�<��7�	^�[�Mt3�f�� ��y���x+<��J��C��jD=��5�xK�R�0��Cz��,�ʟe�Y�MX౨���ڰT��b	g�L�x�.�sj­����ܡ�����f(���l�n�0~ZWh��.���W�'��#rc�S}��g�a׋�)l��|a�x�{Q/����O+����
�ʨO�t.���k7�G/�d����v����=(n�q�lվ���SpO◳\CN�����X����&~36-�`P����E��sY3��k�G"�(�TD�d�OQ⣥�o��}T9�\B�C�``�_��82�^U�p��]']@L�7
k�sI7*�@N~1c#�8�g��(H����ç�]^�y��'���WH�<C��SD�,�y7q��Intn<u>�k�C��4�ګ~S�G�d������Q)-�YA��J��ht�����7�����h�F�Jy���)�x'u���6�	�[m˜����!��;u�+�'LEqP���ݤ1��]{�Ik5}�O��4��
���F+v!�tNQՊ@_���γ#���d�ﵖ٦n3Cӝ����t���!DN=T�_@����B��F��QV� K��g�y�%�ص-�Ȅմ��#��UM,&��c^�`��c���	I��2�$Jh�4u��!HNLR��I����K��.R�����V���y��y�f1x ��{���E'7?p��R��sǠuյ���8�7�Ïڿ`����<,��%n���{J�s��vd&�B��$�{�Z#���[=G�K"e���ר��R(D��9��۔2�,���VF��r�^ק�35�9[x
=O�`ѻ�_+ӰM��I,O��:���+���3���bn�*����= ��Y�U��J\�`l��\Uˢ�s���lKR��7|2��F*G�In~�֣zr} �۵�_�`%�
�ךZsl�<8(x���߬�j�f�I��ǩZ����:��٬~�z���%��v��bb�����6����ѷ^/���>S�}��o���c�Z�ں kMmb��5{)���Եq��<{ӧ:��ZP��$��oí�5@�r� ��K�?����ȓ���"eh�K��(�����.؜^`q��5�*S��}�I��^Lϯ�1�Gq#Ws�� ���(�+�f�1�m���o��]��ъ����6~ANze�L`��z��$Bs�洹�G)�<��9�_ jn�h��Z<��/a�6(d\3�f��a�9�!0�����<��>'���NU`e�i��D QZF�9�D0m%UGc�@�X;`(e?�}�K~|�In���]�X�n�v�@.���Loҋ��
�Y�A�vDG]���m�K��3���HE0��A�ѝ��r|�<%\d�~o�KʗD4�*޴V�~E��a=��J5�@ɊT����yZ��w(3[�W��
�y��\4��Q-9W��7�`4��*��1 ,��} ��r�-EJ�üv��?;�3�|z2�����$���/��W�fk
a�f�ڂ������&�Q�E7[��(�	�y��8!~��Oy�2��L �#�	;8�R-K�U��A�Z������p2�Lhr�U��Ev��@ՠe����\�@����h4��r�;����hϛj�yr����ı��.\�]����]���L
mL׍��8�|,�O�i'9c�s��.�Al�v��n��8�*�����)(���~P�(P��^]���x��LZ	T	��I�$ڤ��hP�9)�J�I���jm�憠��ꮫe��V�1���E� �o��jP�3ȴCK��1G��<�g�ձ�!M!�g��D$o�E{c-�q��:�p�\A�ѫ[�ū2�����gtY��C/ڔL���%�*@��9�@�֖x,x l��"��`B�K�?����Q	�������>ɂ�n�iV��;y�F��/0���Ĵ�Q�Ǩg��
~1ŗ ����`��s�2����-��/�n^�!~̯AB�����i'�\����7��?��Zy*QN��IVd_0;�E�2Q��W:Q�HMd����.�7����z���Ú-Բ�%��)d�{i5��SW�㩴�_��Ҭ^n5�	 �熎�Qgɲ���; �����?v�o��D@oaה'hר6�ۗ�SZ�6A��Ox�S8��=A@�d�z��K�U��<�y�x܌"���D�E6Jarv� H4r�BT�9��'ܼm�����G�''5y�
e�_��PRQ��*�0�&{��&�Ɇ�mh�a���O��hX�>�?`�yT�@آ�A6s�[�q��l}���E��/�T-yOf�%��L��i�u��Z��U	;>�?ڞ����!�=f�>���y�Q�s-3�����wUH6��/ޑx��(��郯`2ɋ&�L6�ߡVbOx�2��1�Z���$ZZ�Z塥W����o�c�<-5��&$���H?5�Э�?�v��w��n���a�Z�z��Q���);����R�^���F�K|�P�6�	�<e��{�!��C�!!���|s���2XH)UqcB0@]��z;YTz��ydi_u��aD����2؆��UI�>���%b����dg�H�s��x�o3��3����h۸[ћ�g&����Ĝ�*#UEZL����b��kZZBŀ!܃��s��w$��Z:{��4�~��9���[�}��n8B_�Q��(��j��k|�~��'# .NI��*).z�0.,��i����7;p
w̌-'\� ����8zD"1�B|Ѐ�a�J�\s���?����F_hr�,�M��AR�p��`Sl���&h���]{ȅ+��/�eb:�
�9�)V��a�9��4JӐ�Q<m�ϭ�h�Qo){yQ�)YIEG�5�"�=�[��gZ7�|���Ӎ|.�d��>���*��}�v��Z�l�Һ�Qu`���0��H�ڃ����T?��$�֢���iL�+�[�W��eZ�Ä������%�6�x(�X��6Q�.��7jRd4$5�H��3A<�s���q�����-��`�fO���萬c��l�V�1K��H����z��-w��j��E�Y�>̮E2ʎ�8���~�C��_M �u�}����p9W~.z!���Œ��6��c����v�Ěu���]'Ԯ��>��86�Ѫjj-���TD0�.�qq�2��x����g��z�o����%�,s��0VS�vo�+�\������*�X4�`��I�����m
���_��HKM���ε��ZSp�k3�N��u�7�/��aQ�E�[� �r��f~��%���o6��	�/�Ҍ��!��bd��H��.�e��d�<�hzƺf��D�۴uL�@�Z�䅺vT���& ���&����w�@p�~���o�y7��\K�S���w�	���J���-V&v�M���oY6�zΚdCR�g���Zb�a�K4�4�-@Q��?�ڮ��ѯ� )J�O<���+@�؄���3˕/`Ra���J2��غ��=�u�nTt^jU\D��\�.��r���Ɗ���=��WZe��~�}�M:��D�3�+^�iëH3���|��Kq�ɉj���Xtj�����¢Raqu����|�Ѩ�w�������������Y�>%b������m�I���y	��f���v��L&k0���tǯ���*�Љ�+�*K<�ҿl��f�����WZ�,f;���)S�E=��_���h1���������ˑ�͚�x�kձ�c�����.�`F��@hA bM<�O8S;�XYNL��{�&�����nT�l�~]��� �d�O���M?ۿ��[f4�,ڇ������L Q��Ȁ-sn+��D��X�}l��rHMK	�_�A@�u�I���� ��60�&�^�cƶ�h�b���R_���tU�˺��y(�.�Y���%�z~���|��lN�"ȡ�+~\�U�ߕ�f!�z��O���$k�+�&��矛?���Ď�Al�����#��f�>�'�����5$Jaw�� N�Ȳ;zL*5�DD>���y`LD��,7ú����\��kh��N,������ω��{|�LF����־�3��k�=�;+�>������4�?N�M���fx���c��N�BP�|(��&{�p5&t��K_��,%�Z��"7h�ޮ���Uw+b(T)I�$��u���N��؝E���� OЗ���T;�Jч�f[�*K쓺��HF�����7��]X�����N���ү��3+t���%'�:��O�'�u��Z��5�����v�����$dt�+C�&Uٿԛ�j�unݫ������k�|Bc�T���|�q��|��f%�7H��E��|PuF��4D�p��/���:&{��V�%@��U�gG���bA��=p�?�Ԯ�m���шMB�kZ�ᴋ��OH��+W<��@ܯ���z�4`l�^�����x2�Ӛ�q�����19�@��D(N�\V�G�o�a��ZҒg$>8�d'Y&��w���m�Y�e��*au�4]��'�RR�R��6�� ���!�%YX�󤣊��6��H��H�|,��ƽ/�R^'Rh��O�"�4�Tr,U����O�0�[9I�st~���kǠ���Ok�h��������uM�I�������M��Q����}��L�+���UN{N��B1W��d��:5��;Ӕ�Ƥ=��e�@�~���?!C�(m�'����}�2����
-��F.���w�4 r��e��N. WC�}���ܞa�����W����Χ��$��]�R�% �*�Z3s�¦Q2;2��8u�e��s��&��hy41�*+^Z``�u7� j�d|���`�]�I]_�w�󲎃 <O��5�*��\��*=I_�N�Nߨ�S�Qr|7:c�C��|X��O�����D����=e. x^�">Dbi�jF���40���hkR����a�p�_��S�6�v �J>��������Z��5�"Rh3-x�i�/^���� ��9�)TB�����q�3-������X�b��G���t`�p��a�Wص��l�"Mŷ�?i��}�@C�y�����\�#�N"���A�7�_�c��B�xh-%��	��u��������FS������Of��NW
0�����~S\�y��R��$�H�N�8���#sKz���J�X�ۑ4�(���F�r,�
NYV� G��Ǧ��Ʀ|E2]�U��ޞZ����n����䟑��#�M�����đN1D��4U��CQ{�)v�j�s	���%�<M!$���o#��5n�AZVZg"�W�v�r�Tnz
��.OŻƠ���w�䁗�ǅ�&������K�t�r�NtL���H���l����9NPԥ˽C���YDb0�\�U��8~IMջS:t�i�Ik~�M:]ny�o\��y�-�@����j�a�Y�ge��������7�)�x���.l�X:6,�q��+�1G1ba=�W�����/5�{������K�.iB���3�(5]j�fjUM=���PV5��������"yt�o��n5���al��5�I�=��jCב��1�F-�I<�o�Z�k�,�?5��kɛ�a\Y0�]@X Ux��d�-9@=�NO3���*��}��8�)�L�9 �؈������E�O��~�)m#�5��?"��Qd0��jJ�U%��g�����:��E�οuA_z���� �D<N���  �r�V}��HX'�lE3�FĈ�'������^[��"}D=����DO�m^JV��A�I�z���Al���.T��{E���{.��aҀ�6P�#���F����B���t!�<PV܆,No:?(>����(��O��&]	^�m	x�t=ػ�L�	.��>h�J$�+�0F���{HF�br�<�'j[�^vӮ�*�\dk�^��?�Ho�c�@��1�y ���c�eMFQ�R����p"���3�b�Y��~��VZb��5�Ƿo�����?��ʮ;�1U��G�EK\�g�g���%�%�c46y�h��	Ԕ̅�!H�e\b��4�>ʰ��_�\t0�Vj�� L�Z��T�a�8�~vi�����6�0�EO�\�Y+q��M�z�4>�N�1c�ý|;V�Oт�<��Mq ��=mW�)[��/h�QjI��Rl�<S����1��yг���X�N-���#��4H��>�y�J�}1��_zt����N���ni/ӡ�H�yH�a�ﱈI�:��G�(�T3FI�]�}��z�Gf�"zw�8�j���Q���zi�*[�װ`�v����P�H��ְ����On��:�5���d(�͐���F��� �����ꠁ���sdk�+Tx�����2�����[-c���b�@��{25W�k-	?Jk�)�@�%������ۑ�J .����������_�f�����SЯ�z]��\�TP&YlwN�`E�0x@�[l�q����E)��q��Yu����϶u��20�r%K��q��������O$�&�"K�9�z���������`�дW�9�����P���A��(�I$���`Ŕ�؎'0;߉���J�#�9�_�O��d�Z����4W���y��LF������S<݋���cE��-��/�TF���R�F�O��S�l��O�2�PJ<f2��%�auƚ݃��L�o�J�wF� �mqe�Rd#�F�D(�;�@�ܿ��<kt�ңVH��z��E��1����>~�)^>+�-�_�n�
_��a�Zц_P Gn�Y���g'X�;�+Nӝ)��K4��κnAf	�l�z�,<<��Q8m�稦�0X�:�V��� ;�Nd����q�)���0����r�8_Ln��U�9��{@���_�����\��
s�W���1�1�9�������?G�!m� �n��z����c�����L-�M$b�:�?N|�&�S\+�V/Iy�%�0�sF�8 �
`�/�X���a�P'+�G�b����8m�#��4{��N4�t��M(j��m�d��rn�|��o��\SyҎ�~�E݌[��;����#���g��]8��0�>�9�f�	�/�"��Mҹc�����M'Cⴡ���>"�q�Me(�n���= ���H@�"S�\G;��,5����'��5�C���?J�ۆ�r��y���my�Ѽ^G�u2�S�1$"��l����=2��)��`���Z�B4��_�u�mJRc9��l��\(jT+��)����^��$7%�c�{ȝaFi��rE���H5˯�!s}%�i,��a��L���-��$ۢ˒���n�a�����`^�!���h���WD�t�Rf�%K��+(|��(b�:�� @ ��m�l�<ꢣ��n�S0ؒ8)MM�f��3}E�����s_L`>�č�%�����O4��D==,��9�"��];;���ٮ�>�tӊh*�����H]9|��]������U��SXZ˵���}������.�M='O�[c.֑�r瀹�&.���蠷Ur�pZXt֧����<����ݝ�,؂oU�m��k)5Ӛ�j�4� ]�7�p1��]�j�a����FZ���jq�wТ��٢Au�a[̔����t�:��xa7iA�+B ����̌�i�,��?��?�,mJ	��1�o׏�E==[�ώ�v��{%~+>;v��}b���P�� -��Svѧㅧ�ǛY{5⥻U�(�x�4u��0���5N��������=���~�Ą�wǩ2�:�G_'[��e"�z�agq��������~K9a/	���Ѓ�7Rs�J^t�`ߤF:��fnﰳ(8.����8V�,���E�F��,{��E<	}:݁l?wph��?�z�B^��͘ن�wh�SKF�.�t7��2�e������r�r�2SZ���Rk�f/�Lv�N�_&����}��v��/�`֨��ױ�d>��t�ܟ_x8��	awюK ��6g��4��#�(aw�����zG*p�e,^U���)�b�_�:����:݌f���aT�T��'�.؃��u��s(�G�!�f��!j(����5���K��qZ�c6���%pl� �������Wo:z9擃�HX��_Rp?pt�:�B�����\-ۚK�Մ�:U��s��Y��B v��A����/%�����{�_d�$�b�	+�f����,i��bD�%T��qk��b{���Z>�(j롋(ݖq=?}E�^]'A$ҩU����n&�Բ�z4{���tE��nV��=�2&O�n�ʶ�%*�чY����P�y�e�;E{%�)YC�_q�;��0��A���^�������5*)`!����.:��,bG$�8��W&vT8)2ȁ�8�)��<l_Zt�2\�;� j�]�����2���l^J�0I�M�*E��u f�F�_��l�����K���Ero\����&Xp�O��PCv����\�c6�Y�5�E��{Z��K�i;K�<�+N�b��t�|$�8��F.3Ѻ6։�;�� I�e�����z�6^���&	�yz`>,�C�|�H~P��Q�?iYDS���̙ٯ@����L�ϗ��Y�5=��7:j���f���c^)��/p��~��BġS4)�m��g^xlQ&v�8�Ħ���d��aH>���>%�m�_ϋp��Uֽ������ 2K�Pȵ��h'~7�75~oGM#� �[��m��t��rd��$�������'���쬙�C��u|;z�&&���̡��Ȃ:�`�7��?`�����ڣ&��]�Ĳ��P�G)n��U`�_0Q &����}Q!=~��1��:RKz���[8���j��{��Y}�Vedܢ�c�a���[T�"��e�K�i�un�j�Z*N��Q�K��J��z�Z0�hס��ڸ��V�b{�"m�� l�"i7zܬ�]���Oǘ|bದ�����(���N� ?�r7W��U�+
����(��|��f��}��}e�1`!@ů�.	�)
��!q#�+�C@Ì ��\���0�Ⅻ c����g���p���$�T�hW/ˌ�+H>��[Js�Ym4��R��3�� CV܅G�+휅��k��y�:���]�<�6	Z<7�~�)���n�v���N������J����Ue Zn��ut��c]�}<=}��7&�
��Ԅ�]h����/W�S��٪m�����(�`��<��vͨ[a�≛i��_9R������;&�k˵�3 c�L��˅`v������'�HU�(��	�f��&b���9�!�5����P�B�7�M�����V�"�L(���p�c�_{p��ucж��WV�|���3I�:`JB�b��Ƒ�q�I�K�i����.���������$?���]��'�_r5lX�VP�}C����~�uR^u%\M��Ɗn�=�'S��w���`�Y#{E��5S}8#�Tv�>n�<{'<Lk��X���:�bq"��3��Bs.ћm2/y���g��1k[���"��R"����q���xV�'%��B���vf��Q��7ol�Vv '���0�9�3�̺Sh(����5�[�u;�W��ǫr���mH���]6��8>����\>|�m��)6M��ʨ;��¥B}���H��ٹ{G.��0��� sU ��J�nA��e)���rVuG�'?A�}Gc�?��b�~Պ#5=��l������pvl�T0+�7��J/���G�L���=ZJ�i#����g8r�Ѷ�;��vX��-�|�|���s�cz��*�SmA�3���{����An�B`�3�,
,X���8%_���I�oN����K���!�g�dQ���
�=c�,�I�H^��9�6�	󮋻�CS�]�⣬�A�5��	�!�6�WZ��j�;T�x���{bm50ꂦ�F��lz��?�@���`�qK�{ȪNIDn��i�'_P;}���@�q��d.L���Y�����eZG����j��g�#�(��r�� ��\�����P�#��$��3 [�(B��c5z=�"��$Kj-��n���V6��������0oM�Ύ`e���*��vT�ٍ�t���L-���u��������o�6�c�v�,iN�q1r����Jc:�;���dX��:xw�y�Bb���Վ�d-0���#�E�x%�y�/�>Vt�|�\ѣ����h]^m�?H=˃�7���<�q�Z$��S��0�HA.�R�m����|�u7��-u�`o ��l�/e5��"�q�T˻����1����nB]\؋w@a'f�;��~�M�ޱgs�i�-����%��|���7�n@�	�S��<��v>�6���|ع��
��� I��p�1J � �5��dj���g��F�;�Z'�X���6z>{.�o�|�ϕ=�A�����'�^帝���p���G�J}pCi��Y�pG]�^����4���dC�t���
[S�e%���w����h	$"����>R f� x�H�XF%�2���7��a�c�G$�썌ݙ��k�\�!�P%�&�]HK;E]��9m�v�lB���{�xs��(|S����9>:���_�\O�jb�M �� %W�):۞��ݸ�%H��\-����^�D�~~�q���G����gK42N����{���p2~�����.٤�ө�o(�I�E*���5T/�=̉���� c��"Š���rI��'	�2��wPt(��1� ���b�l8�a��h���~�Ų�AIi;R[�{J#=�_^ԡ��B�A�}J7~��J���H�jQ��]�rX@�]sk����#�n�}�I�7�L�b5%�vz�����S�3وh Α�;g3���\����W����}y�,3��N{���P�A��J$�6�jA^���m�Ƙ�ZR�z��~9��-`Z�̻3�M���UL�`�����B[��Z̔S��"��s���
9�w��x}h��^��o�I;9�+{���ܑ��R�Eg�|Vm�{EG�F���0} �pO��[�o�Ŭ��,3Ś� Ɍ{&��[xm{�:��i�v�'+�����e����D�^���v9�mq�d�\K�˱�G[l���ɵ��$̉u,��-�"��ՙ�n�:�*�e�;�E+�����E�9��
�J5gTjܓ=}��)��F��z=�V��n� y��ʨ�؊�P�}�H�G���Z	�j��#x�	���nd�x{i ��0}oN����� V�DMojEڏ�_�gL��u"���q��f����>BDI�x�ӧ��ǎ�U�"�>Vy��7f�v7���1r�}��\�lQ�������@O�	9��eB�H)F�7���{�,���DO�J=�R�*�f��
�����;�}YF#���cޭ˻\��ˁ�2M�R�Ӡ�����D�3Q���@΋f�,�ȑ�Е�$���ppE�(�;'��N�k�� P5|��'����$?�c���;��<��GZ����zM���P�Q&��_�� ����Ý�_����D^�s��dG��(��@�JaȞ�/9�Sm�&�\F��E�x8O�^�Җ��lL|�G�i�i��Z��dS�Y7:`���$Զd����Η�Z��U�������a�j��%�w�������DHL2�6���7lS��� �GƏ��	�Ք�����@�o��K+n�)P'��b�r�Y�$tj���r�7*����:'�2@���q⟆��B)���F�����j�:��6�Xw�67x��L:�n�n5���R������ׂ���w橏:���7�D�p�L{V�py��X�9��>�h�^S���[������h��<��mG��s��i��T^e����Z��:�����G5�qu���hL��B8㋤�']�W��eb��<��2������M����hl�/0Q�w��s��� �i�"��$!UUy�V�^��2y��){���b*;�Nُ���P�`��rj
	h�R�A�4-?+m��`������w��1�F����3B����R��b�:`У�+�Q�L��{��+v��E��Thx�[�&Ӽ �(ɄP�X�n������M7�g4R�w���D�;��K�x��u-b&I�0����!��2T�CUU��'-,�%$F���
�|Aqe
����il,7���A�a���r�~�v�&���kڨ^�����z��ʖn�-Zߦ�uPJ���)�Ѷg�d���G�E�u�Z�������b GJ Q����{Gl��K.ʈc̎������X���L��1kK�Br��0S `��%p�֠��3U�����w�4`��FǿK�Vs�F�J�#�����{�/�w�����m�x�< ����X�r8u��M�ȵ"4dgb��&)�O�cY���Emw:�V��xZr�hyf�CH\��?�R��	�a�9\�
]�M�Lh��C����`���
&�Tf*�d�o�Lv]j��S�� (�	�u;��IՊ���~)�b�U����83��ˏ����w����Wc?���T@�Z��.�QN�kj?��M���韕��\�$v{3�^ϡ�����B����y0,��7��V���y���PO=���4	g"o%^Fz�0Z�[��!���ElT�&ª��h=xP����i]=�F3��G��^��V�,��:ܥ�CHh��lB�M����!t�wk��Ŧb��j��G4��@�2 J9��d�$��ٚ��p�/PI�/`&�!���VN++BA�m*J\�	��-^������C4�tb�w:��Ug{Z�����jL�S'h��v�5Ac��]��xf�uj��h�����3@y$�w��f��V��=��E��d���9�����@��LGc.�"o���ݬs�y
o�_:��d���z�	U��^UF�MO��~��̯�)A��}v���Dl�(��<h,���=)�ѳC_�d�`��>�V�-י�r�,��ޞ���*Y& ,����NK��\Jqfo��6�|a[���ggw�7;(V�{v֓��ru�c	r�Q;�wi�,eٿ�x:d�S1�Mz�hxYl�R6!E%�",��./߾���"@��:-,@ /ax��{ɥ˹��J�Ko��nu���)Ύ�V0��d��ZX\�J\)ʎ�-p��"A!�yV�� mͮY;�HI�BQj�P�FQ�X�!cnżסG�y.3g���{����Ѻ��Ak[�R�p������I���k�Y��:��d:���Ŕ]N�Tg£HE�t��u��Q�=�L�~Ǽ>~��y&��p/�T�z9=l�~�T�h ���ɺ��G��˫����R`��i������#��[�!�����.��4�����A��z�Cd2 �Y�GUڣ	�N毊���,�����u+^����T��R�#�qW�/�9�р�F��I���x��Q��ܩOa@��ې��2Z�j��ȫr�B(c�K�B�>�w66��ͯ�΅ e����u����ao��j�Pa3%�c�Ų��j鳙O����1���u_�]Z@L�u4<Nūfa������k�-RV�i!*xL�D�P��?���%BGX���g��V��ٴ
\U��?7c�6�70�rL�9f�b�m	s\�#���j����{s*SoY��L�\��'��@���R�u��,>%��2;�c<�@L� �CZ!��j�5���5U �N7R���g�J����|C͗��/�9��6�t�"M*s����-R��]��C�A��ڊ��g� �r�Ce�uV�=��i�gc\�S)R/m�T\ȿ�m��6K�g�g��ꂧ���<4n}�=�󖨬�Y�a������T���a�E1���O�Jd�N�����*g�����헮��������ea1�� Ī+���j�he+�C�E��H��M���5@eɊf����`7MQd�0q�2������ĕ���/n63^sf����R���<�1}(/ 飻4L
�o�+.(�<B]�,b�p4U�� �#�T�Z���;R�škؘRҢ�l ��䒚T�� w�)�pE�����m1���T9c�v"̹F͎kzr�N�:3�P>ʔ֒���dY�59Y�Vs�C��b�l[5�-�`���q{�w~!�I��f��Ҙ��P,�E�|�[�9�:�;|��y�,M�=!�}Ʒ�{���;Ԍ�{��j�˕N�u)�~G����`����8fQ삘��(�����p㭂���7#V���ڪ�����ĭ����=mdl_��
^���&�E�FLp�UVⳈ>
<�X Q�B8q��\H����H�R$U��@j"��T��cS�u�7zK55�}�LCZ���T{p�Q�tNz��<��Ĥ�5��V�z*���j��B�~��.؅�cpy�X�g��{�m�c��+�m�G`��Cfzԗݡ#����K�� �Dۃ]���٬ F�H����!�H���`�@��ۯB��,��e��
� �W����j���U����b�����(���? jf������~�3>�f<�� g�4�_�^e�с.j�]�ȼ�v��#(/P����T�Ѷ7�	�N��Q���=Z���Er��]%4%��E�湿ء9'p�{Q�څǮt|���v�|�� ��EFl5���m�A7VѥG�zO[��9�%g�Rl�ڵ�Y�^��<*5�6Z��D��%#_���SE������]b*(�\I��#	X
`��|�qT�|;>�}c_ r�26���,�{��V�+�%3�^�(�f�f��G��D��F���{�g�.ç��I���߸�hw��Ay��5inش��ڛ�M�+Zf�lMu$6t2����q�*jY;���;�C�9��Y����C�,^�V`b͒"�F;Rq|��:�&��L_!N_���;�7�V��.�O�D�Z�!<����ݐ;��.��45?���Dd&HC�6���W�7�H���Ku���#[����Rmh�ѩ�
*�=��p9�{��] ���8Ab���ue�Ft�d�tJd���a����	袃�!DXۯ/�}0�m�z��f<����m|�-���DZ��t�2K}�l�f��5�'3	;V��#q�w�z�֎�y������"R$������8X�~_*�R�0���IL�n.NHخ�cj�U�ҫ]�;ݖh�βH	\O �[H��PX�̢7����l4-�r�F��@m�`�N!|lA5&��b�,q�^nxS����^@����7.�8��̓`�O�=�ѲI�ӥm��ҺOb�s����H�Ȇ�6"sQ�Vw�-l�ꀥ"5�t;~dL��t�t9�F����Nvؤ��"�ʵƌl�Ĵ&j̏X�Mƿ����e�+Jw���i|�Q��pt�.=���gbbNJ2��CZ����
~��Md�?��Ե�y@nAuD�� ����A���"�.���M�=��#v���p�6vn]�D�����9�����
o��^���4�Wh��Ǿ\;�sm����'L����������qH�������<�v��ח���E�Y����GZ��e���i����y����3�?ZFm��2���?6.�3����'ug��b	ԟ�?t;b$������w9f+�r)Ψ�P&�X���գ������V��r��8V�CQ�{�%
;(.R�5�N��T-���1x�5z���l!���J���q�c<��ȼYG��� ӻ�Z�p��$O�.�$kb[��2\�Թ@���rP����ǖ֟AAJ�}��8ֿH��YX�0��ø�h&��N;y$���] ����\�@�Cm��y鄷Z��J�v�����X}|8�K��45�����ABwiz|Ľ�k:����,��9���B���JS<��sѦ[�H��a���6�ғ�C-h�<��S��%��sui�4��5�HU�g~0KBDF�Q����˾��8A�p�g�X�������C��\�M��3���\b[.�oŧ�`�ROkN� Xq	}(��  �_-V�{�L��r�`�t$���g0:��o��^ZBy#u��������.��%fb�P=Z*o\�Z4a���N����~ �S6�����.eM�O�$Ě�&����u�"���~;?�Og���KC;9����������kj��
�I��GXc�C�-�И��1W
��"���U�"@(�k��DD8�cj�F�B�%,NE(��6���){ ���f��7C"dh�j���n&�e��Ǻ����'�@bӢK��U�>�l�*�վ*���GR�a�_? �}d>�����y��B:<�Q�t {�+��,��F�2�js)���:·�g��d�<ȱ}σ�<Sn@ �{,GM��/��'�q��!Q�v �Sw����q
��s�8��,R�9�����C֢��#GV�����;J[��{������f�UC3:u��;Ή�?�}f��@օ��'	��L��� �%|�lG [���Z�e,Əɩ�%j�V^���x������ɻE_G��������~�NY�|�*Tܵ��cQ$��{��9�
O�{�� eC6u��eꄁ�0�>y�E=?L&����g��
�%��z�ɳ�"H��-�MH М�ܓQ��^9_X6֯A�(<����4��8B%T�y�}�j��ʄO_�^i�mz��#m�������V��B����m�~9�M�9^_;-d��Kg�Ι쉪F|����}*��䘿,�$�k�f\|�������*C��K�|y:�{(V�] I(X��'L��?����l�l,���N�{ vO
�o���!��}Ƞ�Q wN��`4G04��q��jj죌Wl����<Y�z��7F]��\��wf�q�$"�:ĨQ��Dx���%�E�mJ��	t��V�#�U2

��0��:����RO���VR�a$v�ߊ˽Ĳ��j��5���E�=�������,�俒)�����$V=�!���
��>�Y��,Qy새�����S�j�K��<)���fn��O��]���J�q5l�f�.	;�,A��5�*�6�ԕ���s�x6+G��p�����mo��柺��a:�ΡZ�dJ{ cL(���T��w����E�C���\��3��wǎ�ٍ1 Ţǭ���.'W�ALK�phy��Β���D4��R�OK+g�G�`�i���y��ު����(���5�a"r�{�>t�WG[V�Q]XVE>���YT�|�5��:���ʏ"�3���.��JOK�2sSH�c�c�y�#9�ѭ�jLX��1������1����Ơ��x9jd�5�P��=!�7�a58�rv��ClOZ)��]�~�DJ�������DbГD	��C5"���#¶n)��"M��}Ys�!��!&�H�=�CEв<zF$7�6�6Q!U!s�dɉQ��'�
��XLH�*��۹���K��#˘�3{� ��wߊ�e*̒�a��~d��i�["`�M:e��B�o��׊�w+Ѳ�x��P�:0�ա�Ȅƶ��x��Q���E�]���S��#�T�mV��K�H�W�Ah�R$c,YO���C���r�U9-N���coj�)z>���!�7@�ӕ��+�OS��?��_��J]�Z���Y܊�rN������>�Fm]A�C{g*�  ���z����ˢtR:���l�P�e<6_��L14q�pn]�:BJL��<�it��N ��q���K,ȍR΀	��g3��ɔ�"j6��AB6��~L;���Pm����9��GXuL��F;��`�%�'�(�d'���*����4���Y.N�����^��V=cu�����\7����G�LG�x�S��я�gɌ&UQi��rxm���թl���"ƙYk�x9 ij�&�֤X�O�M�͔P�Ʋ��>�O�Is�DO����JEkA��O=�38���]�P��;Ѷu����J�u'�\����Zr�گ�#{�2�DN�4@�q�E�jI�����%��OY�Oې� �kC�ߩx��4����4.�`���V7��_�h�ڦ��Y>T�^nTh��1�0��8���<�[of����Rҝq�'���q^�d�X�1U���ļ��+������E��0x���|?'�_�GUm��!-A��c>�'B�=ܫl�hN��N5��y�uç�a����~?ßKjN蕗%�X�d������_��9���L�[A�wS�m�n�p��������^���2�iʑ�o�k� �>��������<O�}�-����V\D֡s1ʋ�h�;u�[e��l�t�2��A�1�x E�E�]v5�r�*m�Q:�,�����7?���1C�t�l%����ɥY/��8�bAїL{DC��-ڣ�cz�z��Vs�S��%v�%�)-=bNd��8?��4�������l�crv
�:M�k��4�Y������a�F`L؊�Q�c���
��_�B�=}i�3����� 	��ix=�&����[�	���y�QN�?�Ƭ�D�1� ���Tu`����*���B��ښ��Q����j`+�z����+pꋶa$����]����u"�*����Q0ұ�g� F��������Y]l��Df,�-�×�v2k͐�C���v��?&�W�iȝ:8B�k9x�8�!^ܵ��c�_�U<�}����oe�va�:@��N`xtF�z�P�I�e!eh�����d�CO^Hz�=�:��f�k�{�[xd^(og�1(�G��R�-cG����R�,۔N�]Kn4���a��К]u�9��̣�٘4ECUn�(��R%0��Wn�1�ǀ���n@k_W�<��/v���,��ο���	Fs���I�X��i2�B�4� ��$�Ы+ �%��� 9ƍ�z�gJC��c�1�7z1k��E��Y���^ǌ/��xyjAvR��8[�LgkwU�)tW���ae˜o�M=����X�ĺ�?�M��؝���5��k��~��ǁW����ӏ�D�y�~ua�s����xx�!;��:ʤ�2����st�����B�wz����!�$W�#��Gs	.��Y�R�'Ԫ�oi(r"�c�8V-w�*�gh��m���{y�W�y�M��y��A��8P�長�����#�y�\����J>+n�KN_�D�����e6�#}�:5�C���Q��m�T&��b�݋�Z�x8J��Ry�J)�
������±V8�7'J'+{���{å�:�)�c�6�w_y�z̲Qw7�A��MYS��\��i����-h�aq\2+/T�xc�HF��>��＜���p��)��M������d��)D�ܸC�cG�p�c�?���R����� ��,-dRx�Q[��'���\����ˇrؿә~0��ܯ�26�����SR s���[���Kv[*�*Y;��cN}��=?�>h<�t@*�'
� ���^��1:&#��y.-$\_Y΍�����XO��k�v7��?@x"��q(��{k��W��ώiI���z�	�Ti��K?դ���|W$���c?�e��c��P�g��N��;*�8�Av��#`	�/����YBaE@:�1)K�r
�I���!vp�5�����L�rD<�lP_�V�^ۣ��(�����(���z2γ"ވd��V]k�Cu��e!��180�����MSt��n�`����<�Ni$�X�O���?��v�ђ�	S���As��G;��z�jj�r��t�d��J���R��f�������g�[2�&����"Q��*��뜎�VC�@FB5+�� o��2O`w�t�����_��Q���(N
e�$ׂ�J_1{�O�e{�H�Qr��avr�>���kC�9m���V�����.^�u��f����;�K��`�1�|/����m�<b���T��j���8�L����syK��L�d�E�I�rW?�(0�X2�|���'�撹>������ٕ�lmd�h^sMq36r���y��(�۽K�S ��&c,��p9����;��qM�W�g�Rm	��~��2���b��)8B�a�T��E���(i���P�]�?�p^~N5�.Q�2}������wR:Qk�|��D������O��f��rg�|MS���^�]����fB�
�!X'+>>1js�����Ǥ���f���Pΰ=�|�)��\7+O_�x��#�q��o��d����풀\��H�ϣZ�.����U�A8�Ź�v�����a-��3���G/T�*��j�ZH��g�n*f�(���L?���pגԧ����Ӻ⼡��>XTJ��~WQ�j=$l�HR4:Q����8��g�rR@���8����/�"��a��򋰄�9E�Tk��K�ۅ�6�e4�p�`�xp0W�8��٦1H���(����?T�7I���Fv(�*�7�#1��*�(���̶?�S��{$=|��4$  J�R���E�CY!=Nw\Ok,z�k���pn��R�¦�`Yx��䔛�B�B^�wXIfT�5$���,m�%B���(�&
Z?����.�zEs�ww��d���M�&(6�����
���#)A}��#��+��o*�7��*�/-]|��ҏ^�-S*g2j�6sw��H`��XR�6��w���<3��k���C�
j%��u��3lN<��Y�c�=�]�H����_�r�NX>�Z75i�YG����1,i�$U������֗=����'����q���+h:�myD��"GH���쑉�1� �e��.h��:��^^nO�L�Gv�'���� .ݤ&sQ��R��mr�a��jj�V��.귰m�p��Fg�
:��"�e���
ے!�d���C�4��3%�V��GW���`6�� iS
��Q�2L��r��S߼��B&�j��J�����'��V�{������'��Sc+UP��9��Qo�h͋O�#I? ��=!ۜB^&X�MM.����AP��i
��uhh�w�W�x���N᧸�«mo`hL6���jW&}+C��R����7b���o��!����KV�x[��&��ߟ4����8�|c�V��ISMN�� ��<���[R���@8��]<�{�8"|A�⺜�,I�ԁ��_�ˎ`w^{�F�f2���Ilf����Ӷ �"^�FV��'�M�7���oV�m�{���3<�� ԃ�-~у�6�����S��Ov�e��LW2Ar���0h�&�y�遼�6��1I1�y�3E��s��+�`�j����l+'����`Y/c�e���S�Չ*/�BaV�
R�����(���ŝ*�2MN[b-�����|%�<Ýن�ٯ��_��%IR����;̧��J��g��UwD��$�z8}�c��i$;\{i)������.��s[0l�{���h�F@�p<l�)�1�砢)C^b��@��t�F�]���8h�0�ME������H��Z���po�aJ�H�k�d'"���>�@뽸��*�����,T3DE�7`H�Oa���3y|K��4$�ɪ6R��C���D�<Y<�v>��ߺ6����6XC�Y�ěË!xj=��>īN{}s�1+�士�B!(����X�ߔE���%���x{�Ǒa��q�&&�(Ij�<J���w�7 ���ٖ;Q#�[�#�o�.if�11!�w���7���_�jhp�V)�!n��̞�|rY����A��E7�������A�Ƃ�������X<�$������Ӆra"��C(-7 ��X�M���;?Z��(B���\\�ӟ�~b	��1�sV���\�BB,������@u��?~�ڧ�#t���];:�Ѣ���r���Zw:Je섾5	��iqJ�ؗ�Wزsf}q��i�A�\��<��-ܼ���"5�߮�����z����|`6]����D��,�|��E��r0n'0͇�#�S,��j�H�F�S�c!AP���J���gఠb.o,�^O	A@d��.�����T�S<�k�T�>�_�}�5<[yϾ��`?p�������ح�G�%�/vS��r�k�OkhO��0�Iﳖu`�n�yH~e������R�K��{݉؂����R��Ln�u��y{����k�LJ]���d"��(��]�՗VB��$�5�P�Jj�Lm�'�0�K�j8�U��J��s�[D�n�^s��ϭ��m�
@�OpYĤ��S��;$��B��d��*P��.���ҟ���:Y�|�w�<��$nb��|r�������-�S�P�?&���ե�ٲ�lQ�i���#^d�����%x��'�S³�Ӎg��,>4�*�s�Y�z��pus�@���0���w�5�	k? �DM�m�k�h��t��$}�LBw��������W��ϱM���:x���*�2���A�Y���>�eȅml��Y\�B�̚r��Z��x���N�<$aէv>s��8µ���@�2B$�/�q�c�IXM���_4w;��ۻ:Ei	��=��7Ds�_ڝ�� ��ai��[ڏ�o�٘3�\w@�|��}M�d�͐��jc��`)�ϖy��0	"�4o��J��~땈+!�%�g����I(�:��ۑeg�5P׫yV?�`<9�dD�v��s�q��֬�-���(_9Fg�Df��Bd�^�,�}�z��F�:���]�c�ި74]�����[��~?���9����iv�z�թ�K�H�3=ʼk��[�*H�4}���d�Bʊ�Z���:�F�!�"��ph���ᰁ�֩�I�7W�kH�8�o.��Q�V��4c�}�hK����D��d���΃@�(=c�c�ھ���&ip�Y��N��N��	�ds};tY����%�uk�W�KX2�3�Pgш߹��_�V:��l1��T>�B#��6���(��?��A%�9�B���ѩ0x���w�L���'�1�)0=Hl���33�s��a�j�E՚�A�����H,ZXW,���L�,��
�w'=(�?B�K�I%�;��*�'�X���:E���>�q�e�j����3�6_�`Npn�b��}��;8���M'�'���.�,ۅ6w#�#���#)�P$�������W�<	#�5�J9�8ؕ�)�ڭ�y�X5�Q�h��w~�SG���l� ��?"�"t�5	��N,�WpLݮ2	�)�WFP4O��9�������d�Ʃ��K(:��"�wHVBW�zS�Z��h� ��vt>��$�Hpt����;T&��P�`�?OF��'��yy�d:S�|å�7j��J��YnT���( ��kN�%�A,Ah��pN��%')^�p�G��Ԟ�[?��hETŨ��K0S��B��4GWҝ�v�h�(;�Q���81rL���	�qe2����5�=�� ��@VZă�$��cޜ�?�Jr�K
�keǩ��.+�N:o�;1v�X�������x���(/��Bs�)�.��њ�����1��\�f>���2/�wz�d�C"��:15}�}g�˝��1W��'h7�J$W)�<J[Q��k9��c{���B11,Z��RBV}�Z�YrZ�m%�B[-�$P�l�ZK�0^KY�>�2�O��C�0ф���y>�&����Lt��!���3^ՙ�z��S�t"��Dꮙ��n��Z)���|V<��Dt(�xS%�?�0`|uA�����ُ��d
tp�u9��KCD�RIt�b�����Q� ψ�N�y�Ţ�W�q/(>y���I<&j�nLe�q���Aw�E��>�G�<5<3畫փma�d$�0���H!�B��uO�(��CK� U���C���a3r���9WA�_���B�=���VP��P��)hg�uC�k�F=���5����!�?  �%ȉd�T��L�`D���+�ժ\P��#ήF
9���-~�q��6���۲�2��4�4ψ�q@D~j�M:д�ڬ>�Y+"օ�!R�
�[<ߦ�����h|��>|3�΁A;gֶ9���R!c
,�d��V�G�z"�=�n���1XJ�����+��<%?^�j >zeXab̰}}�>���q�
���A�W�~u��+��&H��,�ӮF���j.�R�ܧ�4t�!s�q����M�Í�S7���NƓ�V�Q��2�0���Բ���"���
�ی}��]��b��߈�Eo�=ů��GR�H�%�QAy�(?I3�Pu��I����#��#!6Ў�Or/�1��#��4K����ꞩ�]���b?s����B}2? �4ݲ4�M�~�>u��!�;J�U����S/[,7q��n�}���vJ3V�v�7w_�N�O��H+&RFr��N�\�Q��L	�V�n��N��La7<GĢ�R{ʐ�jǸa�[�~~�E�S����~Z�񮇫�6�iTs��_�b5>��arm{I�\��ʼy�9�e���B+N���5���h3u3@�я�+�>�����u��+��W�"��:�e��-B���5�6z�1J���-)�����`��C~��.��-m�@E	��F�[X�7�91��;h�jѻU~cWQ���Z�g�[D�jbv��W�;��<8眴/�JP�X���9(�쟣 ��ul�1*��j'tǿ*
ԁą*���D-'gr�GN��w�Π�&z�y?�RBH}�����u�1�;2���t��E�;���5t��-�h�܁+B����{>2D_�x�^C~�s"\�yg6��q{�Bn��?�`idm6]K����	�ט�k/[g�j���*O?��q�;Kqr�CF�zRQ����$���e�����;>��0�v�BUm��i�+�Xpה$`�7~O�<�o���O�8�q�O��BNL�ܰR���}`?��p�*��#Eo�{*���`���IA�Ŕ�g�2�Z����o���Yu��q�?hr���!v�����G���"L@�5%&7\�/5�vQ6�״��ξ�6��/J��~��D��e�b�l���Lu�������/���:���r��}é�: �3��qHQ�p1U~�3v["<�ߍ�wg��8��x�̊�{�IM�\����L'k's�Я�/�Q��Sڡr���2'�u.&p�6�����7;���h�����yg�	js�(�~&ѽn���8�P9=6*��zQ��o��xe"v�	�xqK�Y��s�=���Z.��6d^��!�\4�^x��D�I��R��fH��g����h1#�Y�<Q%A�r�aӟ4_	ʴ�8�k��׿��lyW��w�s3��v�O�.O,���USա��_QK�x��ki<�??e���JSɋ�ҳV��SF1��B����@�J����B7��U��>\0u�Ӽ�[_�%��}��aA��������$�	7���g/��??��S���֖u�&��Ωxu0K
!�G�;�Gl�H��!Ws�hL�zᅧ��<I�ئ���!=C,G	a�	M��s�ÁM| ��E�=�/m����$���@���MM�H�"C¶We.����u��,��=h2/�#��Ɣ��wx��Y>U���b£c&�h6�q5����%)��*PuYb|��uA϶����e�;v�;z�E\�CySg>ac�fɨ��yNuI�D��Dw�6Q������r��v
>� ����#yc���`Z������-O�Ҝ����f�&R	踅���g��d�5O�6��=�E��:"��L�'���uX�[b]�zj�j\[8;����g�U���&Z�.{�9;�~qNSv o��h:�e����>������x��n�q�(��Y��ł�tYf���7kӜ:q�O�|՘8��ȉxEcm�]^ؓdKJ�
%l�;b+O9��,�t1�V�Y�}&���_�� c=b�!|.��Jpa",k�,�DO�)9�L*�- �]�H��ʠ�D_qe���qe��)��"��0����[���>�vO����G:���������]�H� ��G��B�M���ݑ�3U����L�	
�؃���/&E~-6�>�������I��u�h��o���v\���+��ZU�4D�R��h|0�ѣ�;:M�l��@�m��rS:0Ԩ� �t���4���i������� �Pf
K뇭��:ڧO�Nt��yV4���O:����eҥ��I�����r�8����Ը���E��@��e�̇h��K1"��Q���	��`g�	{��*$#��l�����8��S���gh�m��s����I�f���/�p\�0�xlxy�*u܂�A��9H�N��\/������]*Wg:8cL���%�������A�_]� �(�(�8|fP�Aӡ��j��{)�jԐ���_��	H!#i�K{�s*��2���)V�"�d� �<a=�T3����͍�Uޅ�j�A��b|C�N��ش��"i��<-F�2�m��27��e�!���E��{(�0�u�X]?��Rޣ���v-e�	iC��$���ԩ�0gM��5 �����u���=����@o�Q[_�QhP�!&��u?����a����H7���`Kl��aQ�������)�]=��]%�n�`�ٙ��S)\^�M�	͈RQ+���[�Z�"��8�,���Qu ����с+Xl�����Y�H;z ��9�o�eR����lЧ!� ���[q4O����RBtn'Oj����
�х�[���*���[�{���
�=}�����Ir`E�Q�����#*M懺\U��Ӓ�f�v���n��2�")��D�Ȩ~����,'�j��lTNk5l����*���h�/=�<X�P��P�����䦬��P�e��8&�����HmD�$���B��|���jR
�u��yj�am��%�Vr=	$��#�Sju�F��L|z"󮋕<�7rQ`��4}:����4�(@�ؿO�o]�=�[����H��y�P4@����~�h���ar��ٲ��8���p�lS'ތ‫�:�d�?/���/1&�m&���_B�A۬���T�#@�<Y�sށU5?ئI�@�1���7_W��#@jwqi�V}O�crn;*�'=�G�/x*��Q"���>��/�&H?_\�o��qOkJ�S,��m"���	y7��ԕD!:?0�ceQ�_�o��/�Xlo�j���a��y[�RF����ԟ��[�_3}\����^����� ȵ?"t��X������_-��eֆ�D3Z��O>#��S��
�?z�v�����I��Ӻ%�b '��mS�3N�|���K�"���6d��K���.>��p���<��4�	]c�yi��PS�5�����*]�/�m셂��|���m��S��N��!t�E5c�*�r�Om�kT�b�~/1ȟM��v)�O�����$�h	�zR��n��CS<`� �zue��U�.�׷����+�/����[a���]4�ѵ&�m�}[�.���q��$�+��>���N�T$�Eu;���>~P���w�U��څ<�[�(Z���b�ק��޵�M���-�r�����/�GL�v���S���BQ/���iħ����x��7E�8Y�֤3�'��Y���|!�[e�qRtB��i n�Ya��N"��7;{�H��7�or�p�������7Õ���V���}�ou};2h-�WE�";y�ۧ�K����	��v�8E�+B�
Lt8����
�p�@ن�qd˜-�^��g�^��RO��n�8��m��%�F�7�]��]"{׬@���El�SL��Õ��d�*_!����c�0}�x���'1����T��Ru�(��K�U$�2.��khm���W��u]���|-���ܺoQ�\��POw" P����g�,<��C�5�[���Y���46�~WVE��GVC;�G�8����D�0���~uS���� ��M8��iY�&k�W���k�n�JmDQ�t�~"�J* ��
&��g�겵�	�w��1�s�p�`F_���f~�����=S��� ���(/|v��|��O?��� ��_�Ͱ���|��/��!�6��
�I��M��7��^�K1�;��&!pl�{A�-�s�N4�����a�N\=\�B��=�����i�¡Lo��' ��/�b�1��]T��?naD3w�p�ж�\���l{�PlB��ZW��)����>�Yq<�`E�m�fS�Yu<�I*eIr�R@���:��@��->�ɇ����`��
%�����}�ֹ س�,5���af��0C?.�J�t'g� ����l�C�Ƅ�)��Q(e��<?x�2s0�>x���������V9���(_ �-�$�h �`�������5��sf0O�g�!+|0O��[�����@d=�A��p ��
o��@��D�Mʓ�+x��V(����Q�7�6B���OӒ1&v������9��:nv�c�:��#K���@���a��I��N�*Ӗٛ�O�E��L�� u7^�v�9?��7�Y�$g�O���9�$�Edߧ��5��������d0	^��}q�q�mª����8K;q����+��s�ɴ�[*R��Zf�k���Sk�s�R��ͩݝo�_ ��nhڀF 8!�<��)G0�SH�`�?#�#��4I7[��M4o�V櫝���Q>����*'�H(�P��PPҟ1,$\e�@�$^1�[U�����k����C�@\��K�خ�"[�h�\�D�����j�U�1��� N���^����wB��M3
���#���O�ˋ��.X#����9S-�A��q�̤��PO��%��í��70���1~M��{���jW%3�څcA4�b�B������@�Vx�W��E���q"H�������2��qV����	��M��H(�8Q�[�wv��9(��o����m8�3 ��LY?�,DҼ��XWo��e(���O3#:� ��Ц���	����w�F KY{g�:�VEp��L�K-�է��Ũ�0�ܱ��r�����}�@�N�f2�ٳ�T'�ZID�*��?�ɀ��I1�w��;��K󷝈�S|�k��&��� ��iq�<_�i��J�R}�����6�#L�/$���dȾS� �w�7�S[�*� z�E�fsO|-�p$V��4�F�}��K�t45C��YL1�Y!�Z�%k�m� �hN��\L�Jݸ�֧n��%6�,��	�A6`�]Ajg���ᶅ&M�����;�|%��s���P�ݕ�R| ��b�_���[�䎳�Ϸf��dCR.x®n`$ 9%F%f�T��޽u��x�
o%(�!X�G��>��3ao�Q�l� _�,w3��p��7.����.màjx	�~3+6��
�>1��3U�K@�g_�7�r┣��Nэ(���=�U�P_�lEI:9�w��P"8!��z����C8�ED�6 � |���<Y-��Ym�����?�e2yA���l���F����z;H�3�(�3~�O2���Ҏ}��:����q�~{��T�m�BC���H-f�˪�lG���B,y$x�Sj�?p���ۀf"l�ִ7,	q��z>��fyA���p�4Vb&�70�}FV�m/��L��B��B��AqF6זvO�OQ����Ъ�����3���k) }2	1����GO%%٨0�-�S��7͊S1m^���.K��
�޶6�۸��-&���B�Ѡ!��Џ�9!2�Y�`��$��ŭ�t�$��)�)�sw�t�u��i�N]�R*邟���i��!��"��v1iѓ`)0����Iх|3Ք �Z	�:+譩%xh.D�L)�>䖾9ۥ���#6D�k�ϑ��/i&�qngz=K�"�-������0���|��'1�k�D�k�P���[up�Ѽs]�R�ᆸt��}J	�9֌�b�Ùe��ɆU+�7E<,�X���-9�0�~��Za���Z����~_�B_ա�4s-�&7y��!{�ܨwߣF��L���E$D>s�K�8���>�@t�����V��X�v4&�o��6p饼'f UJT=8�Jo	n΃֗��S5�dt��g$�T4�
�f��m�a_�M���ǫ��)��[�K�Oε�0U>3��%��~�ާ�=sQ@�#7٬�%Y`c��� L�M��� O���S�&�Λ��2Ӵ�m��pR<�jsc;nn1 �n�;ACLP�4)��6�Ɓ�!��vt�;�=B�H� ��K���-��:����\@5��%�����/�����L�"/�J������Y&��)]ȗ��o�Izf)���w���Q�n�����b�"r�ؾ W+�_�d�!���FcRT����N�­pD� �C��������t v�u�?,\p�]�m�+��d��/�9i`���r
6��]���h�@���c��V@ڒP�Bվ��qf��x|�p�����~�����7���wO�Z�3�<���L����H�;�+m��I��Ć;�%�PoL�f��k����I�5�ve7�f�-��x)����ۘl�*m�����Y7����_(!���b�\@T.�T�����Y���Ͽ���H�̷�Pk1�V��l�8龒�Ȧ	٤-76�0�pZ�=�h�s��G�t��o!
N�5WI�t��bc��^���P>w����w��W���ű0��8o�eDW!�Y,O��cs;�&�� nkT�y��@�FL��(�v��Gq��=*��|��8;�ǩJ�������~/�]Ls{2_cnzBZ�4n��<X��{��x|�5lb��Q�; o�e��r�-Mnp͏ۓ���F�6���Q�Ź?�G�s����f"q�w�1V�Gb�T[ߐ�/�q�24�٭�0�{J0q�����J��+���U-B��g
ԩ��I��a��,��Y�E{�Y
Cb��7ߔ{׎�jb�ް����t?mSH�z��\������O	"�o�V�G��yd-���g��ܐD��x|W#��jՠc�|���(���a�G���y[�<�T���[]6=��NA@�νb ��SN�]\Oo��(i9�>ԟ⚃�Q�؈��{NB���U����� �?�J�9{�r�=�>뷱S;j]�S����#����{S��rG���s��A���+<�j��	���T���u^�(�(9���$K���t�"]�ߖ
�Z:q""ڹ��% ���ė��}#�!��n��%��"��h�ࡪh�V�v%S"o�п&C�a�T�H�L`�i"�\~�ey4Ux��G���q
�%��K�Ϝh�Q��j#`��(K�~a��6
��洋�'o���
a������{Pu(�h%�B�6�U����y�rU>�jD�^K��-O��ԑ$����[\o�L��Tq��wJ��#���}���e^�t�QW�谰I��I�YK���&U�,Jp7����yXCe�s	켿��[�R�o��M��:�;(�2�ZWB#�Y�Ǎ/Ҧ��8�E R�n�f^S�c����.�-�	ǁ'�N����ŶV��'�f��+-�
79��r�#���Hi�	��e�9a�c�:Z�
qDD�� j�7uf	٪M|E=��[* ��W�E�S	5V�u�S>�G�(��s��ԭ�I~A�j�����I��NN{��B���/K��9@-������$s�]��F���Tß��7A9�=0��?�s����S<"�н>��x`�E[V�>�FQ���p��������P�-��~U�lNt�en%#��bpZ�^��%���F��nMe|2���g{�DЃZm���LBR^��%�㪂��mgz���� a��
k�8]�o���d!��P��k����y��F�Xw�Q�ai�ھ��z�߳B��e���%VZ����xW�3@�wl,	�Yr)��1�8����^4w��z)_6�\�}�]���GH�F����-�;�}1%��)��eZ�����(:��$y���ˉ���U�T�I�?��UN]��� )©56՛����!�0j[��6\s,u%�����&=�"���	^q�u���01١��H�:�H$J��EIxƴ ̀�>�Y������,P��<����") v��o`RJ�9�s�bϲ�K8�zI�pQ���F�Z�V�N�ac��,Gu\�E	gqͲ�%`-�	0WP���0}��9#j�1�p�Ct<�Y#�(�U�Tm�?�^mT1GΓ��rμ�9ѓ�� �S�����W����͞;q�}UZ[����i���i1��\�[�\��˾$>��~&"c��<Qe��'d�a�]��¢r�X�W�G���q�f�Z��rݻ~cA�(��Ţ[wH
v��
�K@����y���	5v���Ǻ$x��$���C��B[	u_KK�p��_Ʌ��S674����/$rBK���?�c�8v���Q�jp6���o�PxԲf��Ȁ6w�_�&��l�}߄!��)��l7��k8�Ʉ)l�#{��1o��aw�Q��u����6?��F��`�0i����Ok�}�5%����)l�g��o��JcLo�"��A�NS��'�_�ރ��i����^����q����
I�Ac�)r���kK~|���� ���nZk
��J���	J$��bjչh?�F���R�Zr�c�ft�.-�7Z� 񟈹�u5!�+�7�Z����������m���Zv6��A�7��`p�%� �.GN$�*����f��\"��n�K9�55��~�/D6����(6n* aam��N��1=c�K;�t�"j�^_kY���)��G���&w�"6.�nQٻ�z*S�W*�M�[e��U����zYNkX��l�Z�Ga��.U�+�}n��ޛE�hȝ�t�0�SM�_"�q��^.�i-�(��_>k����VЀ��ݷT[�#��Y��}��Ƨ��I鷒JMK66z��ǽ_+E�'/����u�~���(b���RL%�l��j��~���ĺ�E�����௒�v�T˯ 9�'��%F�L6E�����ퟹ&`&�H@Ya�Q�b��7��4��(7���g�$�~�.P�����&Z�T�b��ѫ�!Cjs}>���b)-�	�1E�������Ȯ��+�7�S�,
9F���QE�G��d�Gn�_����t�=X26K��D���*\gi�B�A����JD����˞���L��y��[\�L�	[��:wP��y��I���f����b�	�9�����C=�F,f��U����!�]�{z�c��K��7a˻E�&p�s�Xy_#��k��g$q���N�1�L(�@ʿR3���%�b��G¼���M��U��0^+����̩i�}�T�']��|І��m�v�`�~].ܧ�3�co�����U��'"#xm+��Q�v�_����I*��/1S=):M����5�k���������%�	�W.������xИxgD�l��(PF��Ny����u�+b;S�����;�as�t6������-ߒ��S&j�ZP?�U%��� ���D䲸��ηFY����� :�r9;����,-�y8�q��.����Y�`�]뾺Z��.�AW����@B/,�7�k�d��|S#�js|�� M��^�(?�]����so)�k��D=���䥬��E��&Z]�R�j����X7��98�3��ڽZ��̓�C��R��c����͕��c�d�ēE��u��#/�feuv4��n٫�E��$��AW���i�Q���]�����J�K��F)<v��ôR�e���ё��Zऽ}^
*{�h�a>`N�p�\��>��6�7�)�3����>��ckC�kN�
��\	#���24)�md����J����k��%�2j.҂iJ!5&��f��i�m@z�v[P@�$�!]���I�7������]����O�G��~�@���Wu��^&<&�mF�!?�xoF����&n���>"L�T�Γ=�>p����l�8o'Z���_�}m�=n�$�!�?���XO� �S�N9*��_���~���W��6l+l�6���۾���^��b#��)�/�KE�
�cL����tuZ+b��O�:��h��w?`���]Ʊ3a��}L�t��w�+��o�f�(�* 47��%�mQ	%�:%�� ^��M5�N�ٹ������D,���ͬQ_Z�zd�خ�G�<v�$�l��,��J"y�_5����cЮ{��sps#���`x9��3����=��/����p,]!~O���ys5g��٣����aR�0������E~�S�I!�)M�*�dF�r�a�Ņ��< �}��>��	}�k��o9y���]��=!\td��R�3%�A��Ҿ�"�e����z[�g�|�ӛ����!�D,Ѝ�Ii>tB+מ* ���fP �:mx�Skq��^;����e�h��V$*R�+�gT�I��mf���w[� ~��$����xz��L���0?��׍(W��Q
��� ,(Ѣ�%tΌ'zM�%ʓ��O�A���@��hn�i�+�A��Ĩ�7|HPl?��Ur�V�Uz�P��ؖ�~���d� /X��"�b����̓Xo�+�,�(�t��8Jp�]j�-N�p�+ˠ~��U�����^��ϩl��U���ݠ ���w����=���neb�ߎIt�k�زl��Z����� ��LL J��,�մM,���)�,�PX0e����R� �O�C�i����A����\�z����<>}9챙2�Qp��[���M���Ϲ�o�p��J�if�c��p�	�]�F�(QY���EV3P`'�������LL��a�|�*� @30�ͺ�^��m.�=fb��{t
6�1�p�����ms�nY�KG~���ٮq D�0؁�VP�T�+��#�s�)�I��o:�΅	�┚9���fJO�dI�ǫ�qu;���%�wR6X�x��c�`�VquU]��N���ޡ�62����7��i�!&0�b���Rl�Tm��b
s|���$�v�@ogt|,ΰvF0��i!w�O��������|���Y'R����=��2"�W�=������󫱬SVbf���F�R��[%}��}2gFm�P�� �`6�Y@���Ќ3v!V@"���s�p�H�v���O����ܓ����r��[�]�l��@>��MnWk$:"��O&L0sl&]�cu
Y�.*=z)D~ϵ˘t�&��P�X�FA�׺ާt�`LICS��k0���28�m}߹��h����E�r޻T�53x.��-���9X��OY|�ށ&��!��4��MF![��9s��۸���
���	�@|j���f+f_��]��>���x��/�8r�&l��Ǹ��n����zh���$��e?�t�\�-�NJ���1T�L>��utA��j�{�&?������q�v��2�>ŧ�+��Hf;=`#��=�;��z�������rgq �Eb�Շ�p�θ	tv����i��|�= .��b�R��;��0�����1����$A�W|Ƶ��'�������ba4�D�:8�6�_]Eǖ&�?����_jb���\}���P��d�B	�e{iS��5ne³��6b��.�6�=kZ�e�O�=��bVL�Z��_��ds�K���c��o)Nޞ�}��7a�kJp��όP�PN��%+��#*�BM��߆����ڐ�N]A�5��Nڭ*�N��++��3j~h��Y��:Au�c�c��7عq�r
LE��邚��g3�����-R�@�A����6"y��H�x��=�8X�N3?���T�/_�������_-����9k<6 ��t-A�IX���E��a&֨�֝�Q�iQ��8�ͦ�4�2��3G��H=ջ��PzŽ��^��Ļ?E{ #s	��Ԗkc�&5m$U����r��M+T��^.�g���0�S�gu�_�	V����>W�b

w�pM�k$��Xm9�G���Lk㺒u`�P��5��"Oxw]��"5x�Iiqۄf�!3�{�w,r��&)Wy#!����������Wc��-�Q��,!����Șᣖ�Qx�'�ɽ҃u�J���_����fy��D���|^e*�Q'߳�{5�YT�_g%m�/�<9�!�M�ښ5im�>T	*A<F'��Qk���R e[�ԣU/��v����k�"@�b	�N��Z�"���O���� UT>�ȕ�(Ŗ��lX�}�Fu=L,Y�3-���vAe�qjr\�p��˦�gC�IIU@+{a$����t=�L�|qb�^1��ҹy�C.Cӫ�;� ��_��Z6� �?촡�����(�Z���l�=B���>9�V� �l��L��q�bfb=6�11|����r��������0zD��q�2��#�y_�R��@��;,[��k6 }(�jnϹ��:���Qz��G�:�m�R�|Юj_����L�<\�Z�h�;_����Q�h@=�`^�G�FF^n�&�˼�_�	SD�$"�P���ڊnD��x�}ݿ�L_0/�4xԗݧCj��+���ˬċ�
�cp�gF���?�x�Ǻ-���aV��8���?�5Oz�U�m��@1����ۛ��ԚF�&"u>�oq	�Dk@�����0�{i�v�cm.(LX� ��4�aߖ`h�Ѻ��Y,�}E;K���k��|	ʹ�H�8r��C\�N#��lL�׫M-YӢ�8g�48�z?M��eVەr���v*�*X�Z��a�M�-�HR��B�ED�)STT�[$�؅>����8�쬕h���&Z%���*Mҥ�^�8~h�!a���Wt��ҕ����}ϒҜ�ROiu��IJO�t��/5�S�T�޲��)R
*��b>�}��췕����=��Axh����5j� �&��KsNS{#�9�X�szͨ�g�I�d��Q A�D�����I23ϐ��ݐ�c_O�4Iq
r�(A��U�}D��uنC�t)x-���}0B�p�I�H�ֱ��W��O����H����|�S�A�p�f����즎�`��t��.t�5���v�\�(l�@�eK@���%L�<Jdc��73%�
8ci�퀘m^5��`���ˬx^�$���s�/}M�0d�7kɹj>�JÀ�]G������j��?��G�	���n��g��cI�u.Nr�*z7��W������K�ZeJ�{������,�ۂ��[ra�}B<�ķ"�t4��S4c!��D�M���SN�6���)�o��Ħ_���r���@&���>t3��̧P%��ԇ��R��(�Ne(�Y6�Y�*a��37��]DR��PA�7+��S��L��BbVԓB���E������O��:�����F��Z�U��b�X`"�PB��Nyf���w�\E,�7��x����RI�CR6@a%_ T��T��`��\���U�0�~��
�~�$���
��H.oq�����&#fmϦ%7TDJ�MT6%1K�M<�vpV*޺
�I��1�C
�V8u%Ǐ]�ZX���n3d(��{r\ʶ�9�Yӓ�ƎF���CWT�������z�V)���X AQ�Vi�o#�wfD���A'�QoS ���f^�!�HX����ʣ�)�PR~�Վ\HX�Fe�,�S�8u���S���?�6Z�n�C�@īa��r!t�1>5��Fx#�������Q	jhlH�'&�8�푩;O�
̋�g\ ��8�֭�֥�)��
!��
dY�LaC3��mM�6��cI�IA�\����a�>�w}��뱯�U7ݐçP��%�N�c�Q��:��9�)=��)���ƺԕ����	�^V�uqΠ�#��#p����	����詶`��='�}�S��AtC3|�2a6�ADT�-�Z���q�0/Y8�yB�� ukV��dW V�SmVb�x÷�h}2��K<���=��=�>�F?B8��|�� "�O��^��L)�[M���9�|�c�XR]�;�GtA�n`2���r�봳�"$&�+�ɵ��xt+�fsE�����+		ێ6�r��j��bܒΑ"�s��&�=$Δ�ۈUi�Kě`y-���U;�'?Y 4�(�s$/�J���?NM����?p�S~���wvUT����Q�+��8g������:�M��z؄���h���m��}1�-֬��q�����:������i���p.F�6e�84����|���Chj�j���!�A��th�T��oѬZ��|�5*�%á���������z��U�̓b�'@���x��#=�!�In����Ì^��|<�{�B:o6=Ev�WXe��WXes�)�4~�Z��e-��ݪ��`�O�4�_����ZǦu��FD��D�ttL�����Z51�<)*��Q��m�D�!!�,�v ;^�.�U��v.(0��&S�^-B��dg���Ę����٬$�'�Q7���k�&R-I����GY��1� ���v�)B2Q�g*>g� �	pt�4�����S��|���k�Y�ľ�ټ��`+�:��4�3wq����P��J�����D%?�Õ�1�k8E���ޚ�6��b�ve�����z"M�����X�)�j�������[䉫��s�)��q��dAE*�!˗�(���;���"�~�Zѻ���g���'?W��v?��-A�ܨ݈��Ǻ�L��W���66gS���.���˥aR��8�Oz�>�_'N,c��e��q�v2Rk0~B�f�M�xw��A�)��aY�O�?|c�^`<{8�=�&�����g� VL��cJ��K�ŝ=��/fLVCA�,`9D��0vO�&����B��1(;ɟHd���>�lnh�o��y
(!o��j�=�jz���_B_�kS��BA�
��1����#������ ��:�����@��IV�o������Xp��^�@�$2�t�sO�7x���v|z����jq�Ga3XD�C�y
��+��NB�1�P�JX�2l6B��B2؀춤�7v��?�#�R�Bi}���]p���f���i�ٌ2X�gx��=a4ۣO��殛��:0�O��c�U��1;b-t<߹bC`"��<|���ɻ���-���z��Ч�$"���������(R��k�q��i�p����� SA=ɡ���E��7L�;6!w�i�30zó����ʣ�Bz֯�)B2�K�y�0�،�L�:J|d3�����)Y�Bɭ��"�����Ĕ�+v@�r'�%�F[���y��kvӉl60<�5�y�橻�����0�ap/���(��M<�����p��^��x��O��}����Vo��&�[����*�fC#���M�Lr[l�h��Y9VLs��i�5��J�8��
��"^́�>�5V}c�a�V�!��(��A�!�>iܻ��dV�`�����4شY��_� M�����Ǜ��"���O�?lR��p{e��L,g�O�M��������f9dy�v��Z���&��>�l뜱V?Vj|E�I�
L��&:2/����ƌ�2	Kzi��������uV��0�tb�|*a��V���w]kI&/}��ݒ���*��h	
�J:*4�Ļa����y���vXxL���f6��7<˓�.i�zKh)ۖ��,b��r{���3B��/T�zK�H)�ۢ����.����Q���)sz
���F�A��GW�h�:W���X��W�V�1��Tۻ+��=��VW�^�_M�?�仯�ry|�4�N��L+��s'@%G��j������YiB����fSzB�1����D�ɄzߟI�����Y�n+Wle���LM�q~5��ۢ<¯+&2�U,�1�&�}A>
n%�1<;v�v��g��\'w2j��[>�|+�j����0Œ��@qL*y2㛮}�ۙ��n���G����j�E����|�!RJ���ډɄ�)�%|�K���
�H�����~*��J�惒+Zt�	���yYϯZ�b��6��~�ɔ�k�7���iW�~��������e�0\	�	]�/��"=21���;y%����6-sm/�=����1�V
)8�٫.}�s�.�/��b�g��7\�1V�m�Xsc�0�j�����zTQ�D$�`�ɱ�\_j��a�I�cL!��!�2�z�C���ی��a�N6Y�;pH�Z���Of��&�=�E�|���RJ��WM[���nw�T���Y�=�Z�>ǀ�az�#بf���0��Cv�V��m\�\�� +v����zUq���Ϧ�H�؂�S>�~����t0�g�F�tb��4���}�_�#1��� �qB&;��J���^��Q�\��ڑΎk44�4j�b;`��sN��u�9�z-��J�O��D�A9���P���nx9@���w��z�!�tm��8��KT6����t��i�E!�N�LoR>���Ex�k����IC�f��Y��L͚���+�����#'��YDt�+'�Zk��>0FI���Y&�6YE����E�6����暑��\��R���(e�
���!^���e/?�~M���Wa3�l�g��n������@�I}���=?�9B�b�;
(λt�o��?�v�%A�}��2�(r}B�3�/����C ��2M5�H弋�A]�b�,0�1N���u�	��9�.\-���N��:��%�1�^=�-{�UMo��ݣ���a���E���I
!��^u�)�y�`2x�FH���b~�\���#��#�	� JO��<.�|�!`��I��[�7�O����%	��?xn��h��ׂ��2�S^����^H�1�66ϝ b��O��3��P�Uk�1�7��W�r�N�g$��/5m��jz ��l>0��㟑"U�Ͱ�P�]J���t�JA����W�(�c�؇�T�zG ��.�x�G��'m0���j�.[��Rm^m�	6�U�&}{�ӵ���;��n�;�;�h�Jp��"�o���_�Jq�(^ό�ȋGW�S�]��8�^�O$,}lD�=NU���8-��I�LO��#�ѿ�I���l#:缃jH�� ;�Q�ބ�v\&�aJ�=�QW���@7�=&^�Ë�"0�.M�����K�j��c�)�ٔ�m��li����z�"Dׇ��^����Cx���b(��&6..yE��h|s]���zO�f�R��P1fOW�'Aq��Nn�ȯ3���fa3���7�.�8��n6�ӹB�j�7Уu#tI��4N;�P_1_iP�벂�M��m�{�2e�/��u��).��/�|è���/б6nmP�+!����k�W���������Ϊ:��)�5ٻ�ҍ`��̎YV�K䟵�b�&;��.�k~?�3I�����ߐ��r��D�1qE)˖ &����h��k4lݾ@ۣ�,�����t���/�����߰��+����w
�����$�V7��ݥ��0�?_
�V)<87�@;*���F)��\@�~�ѕ��vt��I�p�E�	L�m��몣�6F���e�yI�����t���$rs8�l��6`��enY�s7�ܮWB��a���v��a�S�~iY>�����\"M%%fV!��Nw�bF��*S�`�F�6����;������q������K��<:_8�F�]����5;�|>,��!w���WC��*e<Ώ��.%�1�j�[6Y�O��)b�mk��>�]T��8;G��57
dD�k��h I�"�:S$�?�1������~3�In6J��Կ��V 6i�k�]�����%1D>�{��+�۱���	���^�W�~^5��>��O���.�`��=�J]{��Ƈ���hps`)��^!-A=��I>i[L��e�r�qT��?�ЅMX"���-O[�^�dV��%���!8)���*�qv
Qm��_���@P4�UC\���Rp���G��8�pP �Z��IL9i�5������5��O!͢c`����Z�o!�����$%��I���h�;�I�	��3́s�5�P#xأ�*"0�,/B ��촉�`����Z�ކ��xn��٢���Cg2pa·���.lrYB��֧"��~�V�O�S.�փ��q��M���@^3�K!S�씷2�Ĺ����fP@�_$i�%eR��8��+�O�\)�	݀njT��xDW����D�g�\[`���b�j.�i{�X�=��6�u���|J�U娷�S�ryF5E���> &���X�� 	�����#x-9,5�q���Tǈ������r�D�v�;���t����ϙ�	���qn�
�W6H샩������\�������Ҋ�6k��� ���������oS 	�~�?�;{�݁o����J��An�#t��s��%�&���!��K�;�|t+�N�T��!A���B-�
��N��vI�"=�b$�oŠ���-���`gx)t�$'�Vo���s�Z�z�i2���j�mg�5d�/�񝉷�0��@�"��������H7oGE��A͂����)n�ˢT�?I꧜��Je!��װ���<�;+k]/j����TefҮ�'v���5�F�����DD�+����7��V3rry��z�u��H��39!��)�(?�Ϊ���B��)����$I��	��Ϛt��wg �vs�_��!�*��*b�-ę6�t�X4��}��|W�{��TR��BO+uj?�5b-A��"���Z�j�14�"�N�c�2�@9��=*
���m�̩a�&b�����b�`h�O}�v��z��W������-i<dW� ���o�A9���HV-T���K�J���jy���_�B�No�N"��~ ?R�_�O��p���4�T�J.�(M$�%F+����+QX���Ӵ���y������z��ܕ���'z����O�T�_}����-�D����Yc~{��s*�}���� x�n���nԸ�U��:�Lj�N� z J��{�V7�ˡ���vQi�6d���]y7��<1�w$zK�m6�/수�b_G@����u��w��e�:��a��Y�k;��gM"hd4���p���ٽV~���(?4�}��p��[x�N*�8�n�-�p�o24W"����}P�r(�뽵�gp�"/�_����3�4�;��2p]�"���W(��#Zz
�2�]cn2��t�s�.��,l爋�s򳮯�䛿'��z�v�&w�}���S<�`���}���fL�9�&�2�A]��r�b�OF"#m�g`�\��["-�6f� ܀Q�[���)�^:�@���F�C�Ǻ�ƱpW�,ڭus8S�i(��j�Cc��Ӱ�N�Y���T6U�8[+x@��@�Ӓ�N����t\4w�\,�����`���%$����+��Z ��{���5R���K��N��6Ri_��� s��gS�!y����y&MO֢��,�L�U�O��P�o1��?�>��R���
��7,�6�Vc��RqmSB�OۣL�ǣ��N��bg��Q_ka}7��'Z�T��Ǩ�M �Ը�����@̣�(i:����%����cP�1)���߁�܁j��,/��t/K��+�Ecf�(r�w��d�.���Z���0��[��3:v솞�G��
_n�H���k�$M��s' �̀aB1�p>�~�.�'��@��1�t��*�LdǺw��|T�d�<v=��L�u]��7��I�&B�G�0��%���og��ݰ��e���jY���Ū�}*���Z׼Z=����3�2,���8���i�k�}[���ٗ���k��9t�W���oI�������F�}>7Kd����i'��m���_:O����8���.@l͆'@�i�Sd�� �Y�FȳȬj�<gn��7<۰� i���(p��-���%Z/�ĉ�DXW��$SYF��4�E��B�s6�$S� ��h���4�O�l�]�Y�˃6�$>,G�3uI�27Y�_�)]� z�}1�y�!�(����Z��W.]e�s��Sxv6�֗�et�����<Y ���3Ac�����S�K1Ι������W3x��0B�&^�܍�o�~�+�5�D��r�<� �C���H���zq�߇��	בPʣ����q�^g��Vg��9�������Nv�����v+�@��g��GP{d���n���}tҘ֜��F�����6����}�g�60������.
�l��}H<�`vkk`��zBj��wڡ}�c��$"r�ss��$�W�+�8x�F��X\�+A�@ߞh�k��Q-d�=�m�M��)�(�c�lzo$>�9���ϕ<��P�#�n�q�x���)�R���c� �U F�@"t"0�?�}_Z�eZ�О�����"t�	�o5�ۭ'&�tJ�H|���O���ܨ-��\LDp��A/�P���I��'9�N�)��t1��3��GFmO�?������B�XE��
��VbL����[�J4A�r���n_�Io�Z�@z�����˶�'~���dcc�7��ѵe5�訉�)����9]VԷ�e<�êj/����𽽶�*#G`��`8P�j��4<wig�#�C-�"|��L0]45A:l���?��v�0�G�ؗt��ȗ�L�r�/T>�2���t�� [�����Ag� �9�M�>jS�̏�O���/y�;��G�9���y� ���J+�T�pFh��i54�.�C>ySa��Tn���9���h߭����+�@��^+TĤ7���L�ZҪ�����50 ��>t�.����h�������#dɿ��Ϣ�k��*�{�V^Բ-��CF����� \���o!�1����Ќ�'b��7P ��e�
|UIW)��I?�m(̜��E���~ai���`]��r�*h������i����p8��4QN+� M��;z[���edʆj�\4U�<��.�}�^�=C��k�@I�D<����й�L�D'�Ӊ��.����8Z�T#tє�o�YRk�������;�E�`/��6�ƣ �����Se��_�G����=��s+�g�"�@����`��yѰ�I���͆��j^ь����� !y{��.�'������H�\����G�|��'g�)z�\N"$���!<>!1�
<7����T�W3�;0W}1t)
����
������"n�u���(�Ok��%њ'0Q|5�Wvro,�*��!I�?������İ��F�FsܽpP(��\[S��e����D�|�M�/Uj����:^_V6��/)O+������0��s��oL�CM��"~D�;;����r;MGV��@�7�7Wn3J�~����y������>�⌬�l����O�U�˥���ݙ\�|�8�6?��s[�;��P_�3#�m�
�����M�q�1�'�=��5D0+��6��M�)�׫.�V��^�}ꔸ�drG�M�|y��]��
T*c��fl��@�q�_AGN�vsO�+���2#M��)��^X��6�Nr5K}y@[�M6[�UUٷ����w<�o|mа�� ����^�`$?9�;q�!��: ��b7�>�+] �Hs��)ML�/@��+�(j;�3N��8�H�Uh���Eܣu���%�[h>oB���ȅ%>^�(���\��UB����L�wq;lخ�C[7H��}8���V�&��l�.�	�;7���Uq<���q���ˀ`��rH����
�����q!�e:l3z)!jD�,tҒ��������F��~��u�����Qr~$<DI�!��.��@&3��(�o9(U�в3�D�j����p�Z(Y��=$V���� 838��%��^ًi̓�]�`<%ܽ?3,f	@�L�_{�;|h֧��ٶy�7��O��D]^����w�/ެQ�G�l�_��;zd�h:�oȪ99B��چw�o��g���ˡ���ڤ�H^���X_�R�K~\��0�P�T	h	��;���?�bfv_7����ʁ�]9�jު�*������#��;C��b���>�3(Ȼۇ�ʪf�C�[vO��,�5���'����}>B����y�#m�s����ߜv��ԅl��4&b���*��y6�R�w'h�N},Õ��c	$�͸�����ӧT=%�i��O�1��	�ӣ�Sƥ%W�B"�~2��N��ӮU��pE�4^��*ؓ����3UR�$[����h��~��`���k��պJm
���f���Y{�i��Qʦ7�]K�w-
$]�9�ưCMȬ���z�'��daG=Z�6ٓ9a�'l8��ù���
���04\=�\�q��4/I@��h����o�WCq([ �������_���7E<�%!��5���~f#�o��ct�'+ ��w�݂�IÓMAK�\��vKzo�����E`�j����h޼W y�M8o���_gg�>��}���qS�P�u����]^)�V���l�ڷ,�&2��X��K�wp9����$�% i	
Hx���^��c�G�l����I�gq�fM/�B�@qE��QI6Tw2��8o�L��h��:��.�D.�>W\�H�U���Hv�:}^@�j�X6�S�R�K�N >P��\t����!�G�m� ����T\f���e$Q�Z	_�Vȩ@Oْ�q��jkc/b�5���n�����(��+-w<����ԖH����RTr4��S��x�v��3O@+ѩ���n7V���G���
�/�ю?�9ؒ�/��7����a�j��]��{Y���x��q�'�^��>�7��$�ο����Pڂp�S����Z����B3l߄�4�B0H�u��Y��'��޶�$�1��8�)�]Ի)�����z�-G45�Ј�ݾ�t� ��k�u�?X�D�4# 7������	���q�Z��
Q�2*q1w�bL�)Jw_����:�1o���M��@�4/��Y�5�0;�J���=L�d���p_3�n��$mH�ڳ��cxn��e�_��1�k�9lk����>��J��]&��۱>���H�YvMˁ��;>T�Eη��	s0�/��ԷT�c�ݜO�ҍ����&=��F�Eliq���2��&/�ɫ�hp�u����*��D��`� ���0R��^Uq�#i�#�L�ҡ�'?�7�t	�囔����|��Q��v��2ӊ%hJMey����|�ރ��*w���%��U���˫~ �4�RZ�@��.x�z��1�V�k�L�JRǳ@6��W���-��ݢ��lj�R܍��SH�}�L�z��,�(��YTĜ9�@w��_�c��`tBsW�c�\>@O��J��n�t) �]њ�5󀅵ؾ�����RϪTn�E�֫�3c�¡���XӦ�cm'�(��'��9hb�O��.^�O��Q+���wN�O�h_��[Yr�v����ٕ������n��f��Pӻ�^�~=�A�{z��J����;3�x�"ʝ9�d���F��6ж��U�\��dT~�����(���P�"��7�R}��cHQG�K,�PZ�}G��rMvS��� סe`g5�����`)����g(@��Jz�x/h[͂B��J]na	�-��^	�}r�ҏ�	1�7�}�N���Fw�
L�of�<E*V�#3�^9}�2�k����byΎ�V�z�=���a�g�+#��� [}Nm��7�O����
qFu<諥�q�k1P���I8���I-#���\6��9�i���KU��ibz(H鍤$��%8̩[ˀ��\�?@{�=�I�n�_{�2:�c�0�aB���ح�f<#h���iɀአ��M��-X���F�R�*�WXX�tv&1��q���X��·MQo5Q�;�j�\I��H�hĽ��~��hl!�3�e&�pm�$���M�f��1�:��D�Ee��s����鄉t��t.����~��V����믆3V�t�b�C�I��3�_�w���Y9�T��O�����Z���`�����.�-'#38h�oG��4*�K.Rz�[ѓ�)���Nl�LP*=."M�c�%��5q�A���g�	X�;Mf��h����ZLT�{�i�	�| ��e�h�Gk�!�NO�����!�:G|IC�jK��hčY�;.In4��_��{�Mt��(�g2j�קF��YX�)_:�ʒ倢��t��vHĩ���u/S��'�s��y�Z����k�[�J%3��j[};�
�@���p�;?_���q�oTqe+��JJ�
�J���i� ����P!*Ԣw-]�I�����G���Z~�&�.�[�-����__3���`�ۏ�S#��dr���`�Tf�[�o��m�(.�e~y�N���nK^��}W:]4��@�ŉ6/zs��S��^z�-� 0�uc46O��T'K����,�!���2�d����#GBe�ݳ��m�yg�jq�-�ݺf��I��f%8i^&M�J;�;=8 �W]����E��dnŎ22�;�E��v[���B�jLWg���-�F�Cd�j�ﵘҔ�4v��抽:�6�L�U��u�j�%n�4,�b ���C]A���>�+�T5꼕�Y��+�#��.$<�D�j��K��������!/ny2�# ��Hj��񿦽��|��Ȉ�U�>��:�@o�Cwb,'
>���be�=�Š�'�U�������.�տM���n�B�M�Yi�D<� ���*Ceŕ�����N�Nm#��=�ˁ�P�����/�(�J@�'I�2о�K��.?�lVV`�����F�� �\K3|���y���Q7��^�_䋛�����<Zgq	<��Q[F� G��H�8��Q�v�r�]�+X����/[�c�[0 �L���[���JL)}�i_,M�5�'��s�*(��B$�4�=w����3�$���.3��J�.�񳣄�������1��'��Nn�&��a˙�`� C���WT{�5a03��c��C%d�ܴ!۟H��ԟ"��u��4�%�һg�F}R(]ݫ�0*���\��Z�1?mЍ��;4:y�;%Y����+��� 26�y��%ʢQ�Y6	��_��Z.��x8���m��^��ׁJy0���'[��pb;+�&�ϒ��ߔBĂ���캌�\ʘ��42��z�M�[%Qk��;4^����r���0�X@
�Et�k�5����[@Y,IvAa!���|�GŲ���V��|��n�*���F�M�Z��-���Z�A�9���{�ŝ�'��$ c\���=ֻ�,\̦jN�}��>Y��#��/=��kS�hS9��&m��j�U�G����Ud�̢��r����۪�����0��8[^ ���'<�A�r2 ���r�2�*�,4u�\,W��d�+m�H�"�O�	�_l���~�\�k��M=wT��Q�i�� f�T�U�����d9a���PR�%�>h-�*M:�?t�_H������j�\�@ې{m����/��j<:��K]���>S�%���1,f<�*�KE�oS����dD���g4���ɉZ?b��_����y�Oפ� �c�!C���\��TXN�$�T� [�;�*z��hK���iH���T�{���-6ݴ�s3U糷�X�mTl����F��}��s���a�4AG/Y���&&��uxOx �b�W��p�����R��8\����;�f=p��'��w��:�G{l��g)�K���fjX�*��N~p��	��F�7�MT�$Ĭf��>��`��ۜ���b�o�Z�ڪ+v��jX��hN�Pe.֡KH1�Mq�4N�=�\K��T�WA��Qf�є�Drq�c�#�~Ov$GJl��B�
>PM��xy=��i!"����U��& 2���z�P}"y�+g��6$��)QN&�!�[�S1�x7���+�)��4ӊ�����/O�Mo�d&ZvU�������ѕ�m��b�q�2MZ�Y�q.'���|�u^���}�����Neȩu2�
�1��qb#�e����ɏ 0ӈ/%�>$=Ǝ!��+.U&ɚ�SC?�T� T���4�!� ��F=�@�t19���%��4I��*@���#�)Ha�M_5�0�O��6&ݕ*� [ݧ!t���y�3��Ĉڍ�˜��ـ���*��	����;��0����&*�*
U���aK�aQ�2�a��i���8�X���Ia��Tz���m����_�6�W-�k\z#D���j��V�c��`����g*�O�t��8p%^���k��ҩWaDk�qf3ͮ�Ӹ��#��+�c�2�m,���l�8�4{���M�we��ti�OŻ�?`DJ�w�f�+fP��G�įު���$�y�	[�NA	�8��k���ZV���8�M��m(�i��/�F܆�t����PǺ�޹�@���?g�A���8zD�qL�|	v�c���Li�{���G���&b`n��(�(�u6�>�F�O�Sޗ��&.�ȫH3^�r�>�V����bV��,��%��x��>�����=�Y��PujB�����%��&{x��E�-N�ݖ��{߳rM���-f
yul?Њ����/¡(�\��VS�m�gPR8�5-�#�V�X�2���9��߷^�6���=�k�Cگ�!���?�S*��rɢ�Q4�Lq'��+�_�P�.Დ�.- �Af{I�����60�1����
�<ᄫ��8 ��<�jq��x������+�鞥�U�GnKz;�{��.:xj'K+팖y���'��Nh���d+�&�̧��
6���/!%^�6,�f�Y�8]�?���v�A�����tg�m0$8���C����|�a��IӃ��_�
�D��2A�8�kv��}JT9�|���t�,{�C��?XE�ė]�i���>��q�a�d�~��Q�愚81����_��h���柴m�`@9A��n�; �	���x�3��7�xD�nĥVq"���ÿP�ʍ��܏Pv^�~< ��P���H
C{����W�P�D��,���P��K�G�#,.�5q�
|�s	�ԙ�;�P�i$z������z�x�=4y��sI�ӧ �����������x��ȸ:̆r�������J�b�E���Y��2��C�XA.�c�< O%�k�������Oo�������D����v�X:���J%Ӽv� �C)�;!����`��^~5�l�)�BNQʸ�n|2'��`��	��_ɼ�4�fM�;��5X���Bc�VGѧ�TBv椇򨣎<#��̳�Bij���O>₤�ޡcP�*V��s+e�V��W���z��9�����1�_�Y
���P4�2N�Vl��6Z�E?8C�">�U��ny�I�-�ܵK:/	�\�P�
>l^gj��[�+r�&�Q(�-�ݪ�C<	�]�i��p0�ܓa®i�Ms�b
\�K�-�� �b�Pv�y��W�R���ܲ"x�Xb��T��HB4�gQ�c<#
��&B��ӕ��J�/!b����^����q���{{f[��v�I�NĄ4�1tę�wy�ǂ��00?DL7ٚO��~}.Z���-C���|"�8�Z���p64�J�i_��O����"��6�U��=t��[Y4^�� ��x���KK�>>6�f�0S���MQ��S�[��PH��	�n�G�k��ן�E����},N�KRC�z�̇]=�mX�[)Ɋ�8��kE��i�:� v�HԅVը���u{�j�<��`����"�%b���&+��}�y�jɊ��a�$�z��֠7�ό�O�mir�m_�×��4�gU��A}K��%��$�mW�C�{/�:��G��UK A��:l�����ns�q�9���y%h��J�_aoQ�©��E��mtu�&b9�7<yd�َ��5����U�튯G�i�����Bv�sOl�����W���!�8_`���B���|=�'R�z���d�˥��vJ3��ћ�vt�4���ـS�/O����AD|�����lJ�Q"u~Ή\չ�q��*��a��O��׺ԡB��#�=;�B��<~������N���R�=59�a��&qG�OB8ZOK�?XK���O{�ETH簌p��_�t!�̷�Q���K�ҼE2���j^�c{"�m�\h���Y��U�����|��r����C�G�C����H�L0'�s߶��"�p�,��nyo��"T�u�	ro$�%��F�\���:}�O wH��P9��[�T����7���u�i1]�٬��k�U�_��Q��imQc[�VZ��G��S���z�U�G,���m���M�U��S��Ϳ��@�����ωm.�_��S�;�����}��m%�	�o��=��c
�k8�����#{%���o��w^`rp����wdw�����.�y�ÐY�М./Y2��-�U��^��� tIrʻ�Y����]�ԟ��|��N����V>�g����ݣA#�K������M���8O}�EnLVI�\} s㌩pE�����y��/8w7��c�!}x�S�D�x�@��Z-����U&��q·�:ǚ\OEgޙQ��y*��5��� '�ie�O�?��~Jcy��fKu.s��?�LŃB�$Ӯ��d����ߦ�km���Ӭ������1�f30�Oxj�.��փG��R�ӉU�b�S㏅���&3��z �u�� q�<Y�y'0��`cP[㤐VD9dc���NR��{��"l�)5
�;d#��.���VD�h���Za��z������ݿ�1�cOA�,���5B����X�շ��<K9�*���W�D_�z��*�9	�F����3��SGȞ����H�u�C{f� BY2�&ύAQ'<ge�F�Tp*����%�Ⱦ�1�jZ����c��ds��ޤ�|�3p�� �_��T�X�����|����h�p�iz[u�c���Ӕ��6��W�}��5���?�|�l��m��g[��ьXG�|<��/lv���v�F�"��l#��e6K!�x�@=d Iξ�;}��`���@>�?�_�h�����{�]��<�P��n�����(N<:��c]ƧRFx�#�F��b��t��M�<��-JL� �*7���Gw��/��M%�}���:d�X��%����´�b�j�Wo��"�3ޥ�ƅTc�r��S���3�2�"��ܚ����&��F�6,��c|̰cj�c��!��)q�y�>�O}(H�&����^%�n�Y���褟,b:U+����6�Ӎ�bȨI{�Oф�k���č�ɓ8�%��{!��'���0A����셧;oڂ�'�.nȁ�FP��O�a�/��L"��R!�4���r����3FYP�-_5ѽ�]��Q0W����V�Y�V]~B�o��x��6�z?�܁�dI��p�T���X�#��+��R^z;E9����S�^���HYi<����;W�ٳF^S��kD��+8�
�.��u��*�2����>i�E�<K�����@�)���!�D#r�0ŏ�������ʇ
���)�C%���F9���%��~�O���ZE����Y�m�(ڢ�ɚ%?U�ɼ�q]1���ȂSR�@���%�Գ����6���\L���D=� (�I�%����\���6��#�HZD��Ɨ�ݜ�35X�<q'1O0�xu���{쒦|��T�X�i��}ySW����G�8Ww�W�E�¥M�m���3�B�ȀQ���T4n��^g��tM�B�=as(&�/��Ti���
M7n��îTz�E�W���0�q�����<so�M��'E�kx$���p�]����W�B<��e��hΜ�$n��o�����3^-L������Ivf�5^R�@qyo�������Fݛ���z)6�S����c��oN�Z)�ؘ�bMAh���?��Gє y-&�������Yfb��;Du:}zʍ�l܀Du��s�.��a<�>���Gc�O��'�گW�R-,�A�m��t_Z��<���%��fI�k��9�F9_����O���酨��Bl�[=IJ�;��~�O�6�u�P)te�ВdAY1�+k��OE� ��p�t������d7}w���ڛ�,DZ)�j��������U�~Z_Y�#=�;DOɢ����H�,W"���#n�@�Fk��g����Aq98QQw�7�)��J��$1��	�∐I?� C�%ǘ�|&��"!w�N�^Ƴ�&���#[m4{��>��1�z��5��d2�ʿx����o�r5�����)�\�n1���U%$�-��86<F�8ؤ�t�� �"��q��(}`�Ku�%I^��'��+��y<r��U-F�׍�ߚ�½DP�]%�c�<���!��� ���lO��G���ji6��C�u��A�Ì٠�Y]�G�o�t�\��.ܾ��N_�����7{[��t0��v9��<���@T�P�p�:"<��{`<Abj�����Iؒ���	�a���k4�G��nR�nE��l6�h�u��,w���Y<�}�15�U���pQ�%�m��-P�xE�;�5.[-r,�����Y��y�'b��f�?��)C�Y��*�E����-hRZN��V�#G�(W�ѧ.Y[�w��y����s[������@�gl�J��Kry�N�����VL
�����}Х;��nX0BX�XE8����|�\�pK�C�R50�^�rsjjzcÝ�]�2��8xV5*��_�R����*i�>�;;z �2�v��2�/�?6ɝ�଀?$��]� cZ9��z2��c���R[�6��2�l`1b�Y��e����y��!��������tGu������41RB����^�2Ű����r�f����73�m僉I����/���)}ެ�ف!��!��]'ǹw��	���4��)|M��.K��g�o����3@��H�Sۑ��ZL��(��8�X�Ͼ���Z@�[Se��B^��*�h�ϯ���b����T�8ހ�۹�[�����ef�ħN[�q�Ia,ڨG����p{1�#A� ��J{��hx��L{@Ĵ� 5]����*l�7�jO��磌��fa��h�׍��BC�ϙ��oq��ևH��8�^T-���7�3~ꡏGn�����)��X�bym��h��f4 ~�S��߬��I|-�� 咬��;QIۆ�t/OXl8�uHO�q�3���K.F�8�m��,�_@vA��Ǣ5����ؙJ�v�E�C��Q�s���(L�|����Bhx�Zq�<�c�-�����5nYy��To�к�Dv�>O{�kc,���QʦM����G�N�e�a�C��IE����I;�w�zIqiŊ���ZM� �
]�#�,�緕F��r4m�
��+B	����/R�N6���`c�-�Z��kQ.�NX-v;~�E���.�"*�"X�\�3_>�d^�lX��C(�Bt^�h�V�*�~�NQ�4'�OYv�ʎ�S#s�	iy��_G8�W���� ��R�@E�E�]�!p�D����!f�oiW&���Ro�t}��1V����8�V��Ó������D��$Op�7/���5ŝ)�M���F;п�����C��ǍAL��Xpث�]8�4�7�k�bG΂fٮ,�1�@Yge=y��.I
�}ԝ"�FP\֒����\}v�'�~v�m����n1$����'oت���DU�	�Ӥ�m�*U:|M6.1��`���m��'_B>=��%�h�ږв�	't۾���� ���;���$y]�aO�D�
"WB��f��+���~�,�VŮs"�ȋoL;����p[Dv>ީ�֑�Q���R�>�
��d# �)�P�t��3g0@a�>,�t�-�A�(	ot��E�_�ˏ�ㄎh��;���a�$��@6J�|����u�:oǃ���oǝ���sg�	
��ڠ�1	c�%Ǉ:R�<��+�f�k��yA߸�Z�5��Q��%d���Tח^Ju�s���QqBQ���2ί7'Q7$���*�t�� '�siGnH��.5���)�;H|��>��L�;T+�����z��lu{B�������H���S c�ˁ��"�$�*���*�ړ�(�;��!��FJ��&�9�,���V��� ��S�H6���j�5);B/� �k���@����~�wr����0��2i��_�Ph3��8��(�y8�nB+��u%%N�2<4�� ��N Χ�����D��B���qS�|��@ �Ii!�e����C�B3.��ػ��v��|�,$��B��w:'��ch�w3��G����A�ND��6�"�f��sۖ^nD��GY3�� 3�<���1]Zc�?�K'���I���I�.d�������Za��a
���+�5��lq6*e���Od�	���mu�@�	ێP}P���� ��9�;�}�IC���j��p����,��В�%��F�7���Q�>�� ��І�� _$�ߜ%-�ɧ,5�����?�E���fZ���X
**�]�������Q��n(m����)��*�<^s+����R��p�o��Gp�<��O�l]�g9i~���`��'��$�C �I��_���ԁ�&������sg��H��?�f�\}��h695�ӵb�nJT"�9� ��[r���/]ez����@�%R#��--�@��(J�,��ۓ�>� ����v)k�@۞�6*�wk!A��Ң��g�Z��c=��?�pnJ��o����G��C���At�է�����V����a(���H��Ky.8���>��W�t��
�\��4�W��Y���?������+-�ڰv�ȱ��XƓ˸� �t@�<#R-�e�ʦH(���m'�̰a��$ 8�FWi��#��Ur*˅&��佲y6�\oD���L#��c�t���`ʭeGk����������_<�n����$�o�>����r_������A4���=s�_o���z�̎ `e�p�x({	0�[k�/�wv���<H��?����nVݛ~�!6���F���/����7v��"�� �i�+TQ�X"�M�|�O��
��)�ҧ��@�_��KjvH�1/���!ky���a�̂Z~|��y�o��n��E� �/��'&A`�� �%-�%�Rޮ��8m��92�t9z{�
,��|����BH�w��ُiY����O��.�ٜ;{dp)j��uNtU��
��)�|^�9��
K��#=�h��!l-NB��7���#F�1�Asy����N�xN\��h�a8���*�l^�]W:��JR�� %���vX�'�{V_c�n6m �F�1f2>|t�����v��C湼�̎���/���ˢL�,FE�Zqj��1lF]�pG��D��W�Js�)��O������;"�8�+"鯄�_+��֎E�4��qԌ�M���7�9��q���ś-V�*��΂hP��T-��D{�����x1��*XB4Vm6/�J�w��� }N�{Z�2�Fo��̜��2�+��'�d��<x�:�9�&�C/�~})?��/�o9��Η��j ��+�s֢���S�RW��-�D�i���R�%�ra>8^���R(5(�ץ��.�-���n?ߏZ�h�mı�M����+P��1"���h
���ޣuS���������VlIM���sn���+�'�����dl�?f���Uv�}�Gj*�����yyRo�G{]Q,(��_<)5-�캾�A�L��J۝�'��~��%�� ?E��E\�5�/��n`6�ޑ�Ǐ��c����4a]�1�l=

k9C�v]�g1�!�#�e�]jO»��' n�T��k�9 X_��*+.���w��˻;BՊ�Wr&�"I������m�MH�+?f�\�ȼ��"�e�vx}�$~��g%��'BY�̏C�8�.�q5��yb�i�O�~.b*�W�D�uJ�uP��Yޠ"�5� �Chi� S�2~��s����8��a_v�����'��P�*��!�p�͛z�P�E�:���ၧOC̴4��F>�4�H��]������/��y�W���DN�7|iƆ��M������Q-�m�Ң����B8$*�&���;�V�r���Ы�_�'���,x1G+�G|��w�7T��_4��v�z���vDM��'p�+�+5����L��MEGodJ�s�"G�?�n��,;6� >U�:�%u�

תS�!T:a�V��r��/���`���<��u�����c��N�R�R�-�LFZ
�Eg��>/�k�FQ��s�Q��F�7G�8C��UcόL%:��aP"� 3�{J�ɷ�{�z1ӥ��W1�;�D���\������J�:���m��`i2űf���Ѻ�6��,�)�pl������$�Ǳ5�&��Pm6��Nk��x�>�l�Oc>� �`�:�y|B�$P�a#��n�S3:��8D�}�����e3J��?*B��xDO�6u����5�l��_k�T�����QL�R�`�F�f�L���Ed�71�m!���u���-�M�,�g5B�hq"����|aY+�b�U=��s�{b��w��tl	E
/�o�hO��󞣳�sL
@�zf���eP�ؙ�j+��ņ�ǭ5��9�{r���������&�}T�g��,f��p�k��������\h���Yr���Đx���ѫ��)�L ��ob�KPA�7r��YK� �H�~列�Z�CFA�'䛽�硢a黌�� a��euM�iX�%=�)��,��}t����MUw��#�{�^i�(fA���N�-*���2��������$	�p�KE��{@�<`d(o��9�<d��2�OC|���#��
���*�;�;����Ц@�ƨ{�vP'i���_:X�>gd�h����7r��J�Iɍ7,t����< m��9HI�WR���`n�ЛՖGe�a:Wm�mz�a�9_��q�s����B�,�Ai���雙��	*��#��x��pI��w� �����p4����jdU�m. ��Ë����6�H�F}_��ō�l�3!HP�Frn7��7d�:���ce��&H�R&�{'|��:���D_�PNXj�gUƺ��%>�w<��;ԃ���ϲD�YI]o`�Jwe���4�X=&9����C�/G���
����o�R�S�
��ZjF3�W���� ��/ӑ��á�Y�
E0�����k6FÊ�R9Q�~�&Kș �m��,OG$u��̩'���z�	=�v\��
F���h���s7;�@l�S�`X����bI�I�� 1p^�x-oMT�$c����)<���� H�K�/�1����syH���&/����-sb�<H���VJ�eat�b#rn��L�`�;7�:q��8M�(�/�T(fS�O�M����CZ��k�we�-��˅��L�K�A�%,4=�pI1�Jd ���cI#�mqRW-���j�z"��q'3;ّ�G/�mv
��4\l��o^�����N�A�P�>�4���7w͠(�$m3�W5�M3��߇�}�e�6[0�f]��}�[E!��w [c��$+F*[�9|���ȹ�l�S�@ⶹ��I'V�ߌ9Q��/�b��k���<�.�B�5OW�M��J;�G;�G�$|ܵ�-�lt�N�k�(=Iy���J�'��4�wX���A���#ڠQ��]wZ�����6�w��Lu�K�d���'�zL��2�+�T�S h��d+k!0��d�A�p�m��z�m���Ԍ�a&(���8�c���ܮ����ꃣ��;u�Q�$UZ[̚��~G��@Y��B�7ծ�� 8ߪ��.)�$�})T�q��v�rU�������Z�-h8���R��cy�Z��Q0��i���Uj�1h����B���[W��4�<U� j�/.ޫZ��Dh�s��H9��ݫR�Eކ�^��>H3�m���@����A�TqUZ6����I�6���K���/ 	�lz��k��@o���!���U/s�ßP�_
:�v��_���>��xk��"E�n�XN(Xaa��g�~U^#���*�b>O��މ��ΚۻK���!w,G��S�t�u`$bW1ɓ�(�g$�N����u*��WWۭ���#��~F�3oM��).�,<�q�=�QƋ�S�o�=�>
���k^}q���������w��B[��:5�z�{�b���v<���t,B�{���j;t�,�y�����&���$�U�ŗy?�*��%��~4����a�|�	=j3pEi.ӪM��{�2:2]��4೅4���"��)��˱@�F<����Pr�U��v�/y��G�����/�7o-�v�9M�z�/�K?湕R?N(au�'����(��N.�^D����7kW���vq\�-c��&�_�S>P[�p2|���H���xy��n<����\5đ�`��g�AU̐Qx�lYK�p�yw�ka��I�C��/�7+�`��"�=��R\z������$m*��N��ů����c���1 qN�=��]�rd�k���0)5+]�?��3��8���+њ��rO61\�B�oXG��KXӑ���<��x2��˽�ұ�R$�F��E���x��N�L?>�0�m��a�^�iy������]\�'܅�D��'����Й㈚�K��i<��,�7�%�Q��Be�U��G�t������Vؔ�"�Dq���VR�]9Z��D��7�X�ɷzx�:}A0��7#��a6[J��j�Im a���y���}��bU<��T����
��+�&[nj�}�;���+��_��9�IP#�H(���Ϋ��ӕ��}���$Q�$^#A��%�#~B���i�g�2��$H9�Sp������.�!�����@�y,-�8����.-)�]��Rb� {8�����D��0�^5h��]��H�_�x�ϕ��.z4�NA��F'�6�$@��eDbvL�\n��r�Q�{�z2HYu�ħ$����t�Xցf���9���2�~�N�v"�v�gx�v�4��PZ)C�u_fam[�PFҹZ��<����%�	Q4a!�C1R��;[}w��`d(��"d'X�P=� z�dR�U�Yg��~����~i���7V_��"�wr��J���)�e*��qz���e�ܡ�g^ Ԟ�*1�0������uW�~m� hK7q��Y��z�D"=O	ߵk�L����s��]����o6?�|�q�v�$D�����}��H�+�iv{����0�� /��s�!�:��(:D�����t�A}������g���
����c�l���r��dZO�W��Ԣ%�n��T�+7��w����b���g����f�v`_�%��vh%�`z]'.
z	{wP����1u5N�<Y��6m�ޟ����HX?�0c�1ߦ��YP��}��x"M�*�+�ޭ�i�?���X�OBt�$4/4KG˟N�˗\�'A˝��t��� L��R]w����SǦव>�����:]d+�CկG�
{0;�����H�c�,�D7.�W��?���HED ]~!�9;��)J���@\�y	�qH�|�
C
�A��!�q�L~�p˪F@�h���"9K�D̖)���!���۟B��O��ϻ����[ļ�-MRv�xnM�����P��Y�R}��U�-���AK���͠c(.��r�.s���1^��x���଺�@Oؤ�{2��,Z��q*�
�t!�p��G|Fe�O"�����'����$]�n��ʃO�l���J��'b�x�մ����d�� p|$a�>��0�gP"¤Jƿيm�RV�a�F�RòO`M�CiLfe+H�#�r�NM߻�U���,o����P�#�z�9��qp���2gjRz���W�ٓ���Mm+��	���F��2~�C��ǚ"�S��^8$��r��(�v��f%h Q����P�.��b�`��k�����k�ّ��xO]K����0�" Ju��3?G_����â��k��F�&[��J7 hhR!��w-$߈s�����x�>>6��2���}�Ȱ��Ԛ��ێ�f�w��A��j��~�1�C����q�E0<Zj^���ݑ��6���'�ak�G𱡶������}>��6�4\��Om+;�X�<�<�ĎKe�g+I����������T�U�n�p<+?L����:z���Oⲳ�m���a����o��B|�R���<X�g�dl�R%O�2�Q��9J�B���TJ�x��҇X���C��7X��5�p*�ݩ3����o��)���:��.%��8�Eԟe�h:�ë��U��
�㱷�`�=J�mĴ������ο��4>'9�u>��l�ho���quJ�<u<C1��)J�1'��!-�f���0oc_��z����YF����XhW�V�|�یF޼J:�Lv��FC"3tϊC=�h��x�=�n��C�C���k��޳B��bv��U?<j�Y�h�{��~�t�+�!T�m�3D�s����hUG������ş}�ժ��;I6>��D�bLpI�m��k	^�H��H'��EpV��\G � N^�y�\�+�j ����/@	 �%�'�Hg.M�Z���w*�Fm%S%C�Wk���
Oa@J��hug��t�f��t�������xu���B�%�9�O��\K��Y��,��O9	��<K�P+���z��,���h����r���zf$��9�f���D����N�(�M:KE�o���ǅp2`e��h��+�趋�I���9(��1�G7~
'.t�Y*���'ɶ #]��В ѳ���0��dK'���{!9	
g���*�`4RU"���F{p�|�0~��1r�wjR��^{+�g�^��?+_c������*?��'wj�Ig��� ��|����:�Xi�N+ǐ'=�R4?q�+<��'�̐w�,�9ө�1犙�c���^���S��zM/��ܙ�e7��<h�����X{�%��i��]�*Ǳ�@G\R�p״go��`/�� �\�.7]F?I��p��%p��j9�� ]W�k=sKk�W��,6���U%%	�F��ҕ�� �]cA"Kа�*��Bn~�t���c���;u��)������vђ� '}	��I��q���'�M����5�_�!4�ܘ��%v~j̀!�����%��{�؃�����t`�0'Rxԩ�w�n���%f1��+15�(��a(_
��8F�y<t�݂]Q�7��&C����W:b��?Y�1 ��>�>�[�G~�V]E��G�5ii�T�����G(�5�X�_�!�vHJ2]"�H�ao�W����?B^u+�/; �O3GA�bM�n�P���(����>�N����;���ؐw+{�m]��#�i܁�<p�����t&T���MlMA�q)3hu�~u����l��7-+(���"��\�lJ/�0��z�ߚe�|���o3=��Pu/�P�X��@�p(���=;���9O@3ʕ�=1�؟w�X�Ϊb���6/���M$	/����»L�]�=�by��$Ta���>$�%
})���j�g�JkFgUN?-�@	�9=م��{F��DG��bŦOZ�%[3��a���t�t!�[6���{�O��"L���5�ŧ��yK�4gT��G!L�}���RI�zmbY����"
�|�OE���P��r^���������-v����3�"]|���2��'G��#�v,X#9�t�C[b5c����Wo�R�н�hH���H(���$$�9��f�wh���}�Ā��P�)�(<�}m��إ$�3�VԎ��N�ݯ�
t��W��u �nN�?'��lE���/G�r	I��� U�?�&�2aP�U��Ņ��$Ƴ�yeq�)�2s�d���)�C�W�g.�N��K}DC�tƅNS���i���sa�0�:�'���՜X��]lE!B�1��1�;��N��U{&B���]'��z� R4�}9�޷�c�SΊ>�&���0L9Ȑ��_p�Q��Q�OS0����b�*�:�d.���M�,��Czl�[��9s��l}�3�ma�Pz�1���y���fJ�G79<��y\��|�X�s-���.��u���"2	
s,�z����X���im����)k�ZK�čMk?w�L����~S�.bڪ:t���pơ8�^�/�X���l"Q��l���z�5\O:�8�3�,����a�<� sc����0��Q-�m���ݱzxA�wR��=X�ᫌ۳|C����W�A� �l�;,�w��3w�J��2��� u��R@�<x���	�vG�q�$����0{�������eB���>},|	w��ޚ5bDƤb1�R�w���gP�dh+�	���=ɮ�������#�%O1f^�@Y�V�
��_r'�Yՠ�n>Ξ�-w���1�x�y����ٞ�����Σ�d��#r3��o��H�<�0�A�Ds�$��dzC�8�9�R�C�lY"qmSm�r�8A$$�v~�v���卬���Md@ �(��m�VL���.I+<�_0Ͼbf���@S�d�J�#6/m�|��،.]�M��"<�������d���1�caHoQ�?ϗ>���lb�B<�T�u]���cW���=d�T����ey)E�m�T�YY������D�H�y�%��҆?d�C6r���M)?$S�u��4��O2DN�Xk��A�$6u��fk��x��Y�~�K�s}�:awE�`�H�ˮv�M��V
�����W2mK�L��=@�/�[Qɍ+���>n�K��~' �P6�kx���_��W��t��\{5��)��{��~�l?� �Ň�ư��� ُ���z,�a����3�.���Ys��*o�L{7��i��F �Aa%h.2W�O�L9�:�o]{c3~aVeGc�-河h΅����1�B��kpWw�\�ix�or��r�EY �ʳ$���o���֑W��ŧ31A�n"~p�TM�x$���
���³&�C}�ѨO�4��q�9M��=ْ�� ��V�ߨ˱�Q�6��/�f�4{���.���7\��q\�~��t�SO��<}�;���8.��w�+(c4�u����d.��fQ���	|v`73AG$zS4�>��CX��1�}��,�&�a
�g_��Q�!R5u2J�􆴋WK��L_Ś3�݅&��bQ&'���cb��G�kd�?@Y�F�ڑ��ٍh=��۫W_8��/���|A4G�.�>�7��"�#����0!2~��i]�	���榔�U,-�+���dc���ρ3����D*R���h�s�pu��,^a�3q�I� AGȎ>���R�Є_׭�I? Ƿ�~�)�'�EA���nv�A����a`+8'lTZ����B"',�aɝ�UH��(�{0HK,��jk�!<�Q�x�������F��&���(�������|��T�eV��6�B������������:���u���x.�\X���Pwzo��<�����X]���WH�o�����@�(8J�8��e�-���^p�+wq���Q�h���y3|��{��%��$�f�D��rt�ET�����K�/�R��B����>��T	k�|�p̃��lE岰?�i��Q��ě�Zz�	����OQ1b��$��<���L����x���Sd텙��x�5�6q�>»F!����,��_��C�������':�|%�g��*4�k)
�=(�6m"�c}N�}k�"�̹�W�;�c����>�( �-�5�Yw���j���w�
eTƊ9�����F�S(�<�ޢ�d�S"S��f���vk���S蟸��C`�����5,���6�C;zוs7�CH�Xm�՘�܀=WTp+����^�i�V@�gh�r0U�k%W���p��{ya�4�,� :U���b�> (���9NbZ���|/+Ƿ���h\;R�E������s=f�O�v�Ţ�����>���!�e�Q�S^FW�Y��.�̿ݤ���/s�p�{G9����J�la�����V�)���t����X��1wr��m'�6$�m-�p>nS�t7z�G,���xx��_����A�I�hu����3LŜ��&_��85�Ӂ賋��k���4Q�"�f���s��Y��aA?��Q{�غ˟�Id�T�"F"a@���H����W4��������*5n�T9RsX�%��[��0!����A{En�����S���UI��B�HXB�!�g����*�J�����NW�dd�"�`ɮL�C/:�i��ر���_��ʐ�=໩IG��qH����cJ��T�Ņrҡ9�C]I���Х�+�x�'��5�\݇�(x쒴eR��o`����J�`�AG��w����l�ifI�w�955 ��Sұ�����ż�|5�u��B�.RS(����T�\�ƩO��"�m.�3�'��
E�E��$��bi|��M���oN7���3��Te&K��"5f��y��KH,wD���w���.�x���*AN#%΅Tx���4=�*�<c�!��҂;.�8o���Y��7@ʊ�L�����M��	J�|A��X=�G �f.�(��\����j�η�������~����$���WRsAH�k2���D���X�n%�T���@Z�͛��A�����Ct*��F�ze����W����k�fIz�Q�y�X�1|��Vg���߫����aq ��i
]����J)֭�Q�E�'��Mj�d��R	]���,�5��gE������� ,�����j&���&C�+�l2��n�89E+��i��>�Tp��A��HT��� �t���,����I׉���4����e�R/���1|�d����`�+�%�M1�����&�z��aW����fp��X.�jg�>��O5��8,�M�/Чr1�^YV�l��@e���*�
r	�&G���x��]R�TJ�g!����)"\/���5�L}�'HUk�	�s�J���+�6�=B�(�S;��3����d��G�l�h"ϙ��ع�[�ZG�	-t/Oy0�]̀@�ԑ���õ��n8�X+D}b4������� ��k`�y�u�v� �lQ��ەE�VEt}�M��OF�)� a7�CS���&�}ʵ|b@���"��A�5(L�V-ZY�4����?4"D����ܓ�>4s8�&WϒQI'��פ��Z(���F��\6ڳ��72r�ayn�3�+�n&|�@6�xB�K�8"�~8 ˞��L,�z����'�M��P'N?���5C�eh�f�K�x�G�����<�Zk_աO>����e�~��S�z� ��'xz���'�1KVW��Gmѹ�OO��O�'uZg���g-#�g)�~�{ă?�ϳq�P!/3��e�&A���w:����z��3t� ���� ǹ1.�PH��\ƱV���O�������O~M�Hܳr��Z�if���T�;7:�T��G�����&E
j�E�JJ�.R�nN���cq�	+�9%�4+�%IZ?;"���G�aZO����7�w��������ꭧI���h��ߴP�hf6���_zV@�A~�m�O���6F�X�vPZ�����'IGe�M��roGS�`u�������Gg)���A �`�)c$���̿0D�@x��A�BpiG=�h��Ձ�g,��f{{��Ls`�p=��@o��?�\M����^O�k�3ћ�?T�qѱ��?����橿F��e�2��?�I��p5���*v�p��P�Eu[�K��^t�����z�ץ>}�d'%}����,�6@��/��שn���Mo!��D�^�ꦝ���Ǘ�����z`�%〜��>����u�~V!��y$z��|f$�T����!���b��D�af��k�G\�C���Wã������mU2�d?��n����j�C�\��A�K)�*�i�㞼^*,'���y��*�Q$J�%{j�~��UQ�I��Vo��M�4T�����h?���E%�������&��ngvM��D��DLKò8Y1&�M(��J���7��l�|}dt��Ń�Ffxy���S�m��2�^��}�Z֭]\��)��Žtd�o��t���UY�(:j�9l*_�l�s�K���7iI7�{���Dxp����Z��Rf=�j�͊]� �h�e˰��&�8r+�6�dFF��"2a*�����T����(j��p_+��Æ��2��f�����y&���R�Lk�	���g5��Xҝ��� �wG.��)���==�'\�h�q��l�Z]�}ZU��P����_r�l}Y��A��G͋��'ݑ��0��v9į���'�:4?6I�-���^���ȵ"{y���Vz���}����/�I0pj��	ݓm&B��z�%�*V��os[ z�PZ��d)1J�r��x}fȅ��qߓF���Z����,R��֡��)���kO�m;:A���)��,�'8S8�W=�G�g�d�QSN�G�=䓰��w�H�p�?�Z;U�6�����C�W|�^���j���L#5�w��t�e���s��h9E*c�b|�M�K
��BG7�AyZ��
 -�4���8���7���݀���p�`C�+1\h�ۈ^��_�Ff��Ky������]tq�~3Ѫ��K�I6��Q��ʱF�,�bp�Ģ#��u�����%�����74�.9Nm��<�A�e�$JP��5H��:��c�A�AG��̉�.3 1����|*��銫>o.��DP�֫g�]O̦���~���*�J�c�n�	��YY�u�> ��z��?��ߢ0/SU�Sʀ�Lq`���,G��<l2^���������}Ӊ͙{���Ő~^@g�Kdѭ8v��҆�=D3�#�M\s� ���R%�1U-w[w�E�a6�e�U1�V���F6�u�%i1�:�½⣲��%-���d�S�N�P#�p_�xdS���LY!��w#$d&�Xw����n�L	��b_��M-�������	�eZ<�?�S�+�9�����?G��?�?xt��D����*�i̕���}hP�G	�(�ˌ*��=D�Q�8�߃c�N�:cRq{�Ș��{�h�h�oPC�����)��	b������R(#a�G�BX67曤0��S�O�U�NO�\��f6��nǊ��.��mW�wM�O��a���*M�i&QsT21���*
��8� �k�ڼG�<�ܝ��\���9}�|B<t�Ƕ#�bx�'�N�1cYo��2Y�U��'�F�C2�k�y�R�j���V4R�iڜ+w+@}z��t��_5d�׌� ����ؽU�E�_��s�s�ā�׈�[�9�5�]�tv��%jp�cC�Tnr�NO	ax���.��'D��A'`�6����!��4��H�s_)L:w5Ȥ�� PR\�>%��3y(F^}(Kel%W?������,�ś�N���O(�<�*���	}��ڳI�)��<=����B�sbۂeO�$J�Dh�n�F߽TA�-�}����j��:
�������ۿ�*ǡ�T� /�-�u�R���`�j���h@�SÇѐ�WR�1'6i��q<�A��о�Q}�?ݐ��r�R�3l�o��M䘔f�:��?'i�v1*cKb�aT"C%���V�� ���4�\��p�r'�Ա����h	D���Wx҉�>��u]�c��8_�D&��.ii��r�i��]�Z��<��FhL�����"����7��`�dD��Φ�"(�}Ijf����Q���D��}$��Z���TC�"Qil�wvcv�&����a��2'��Ԋ�c��>p=I�~�l�T٦+!��iv�ij�BN� [˾�30L�I�k�Ї�Y�X;6'��"�{�Yݒh�ӓip��"��m.'�t�@"0MK��7���=_MH�[D�7{���SZ���F�,&��n�W�͗�e��	.���t,g�}P�kA#�G�H���PL��+�H_4ޘ���*����"D�D��l�!P���?�4�����V���dw��uɄ�76��(��kt���*�LkR�{�Z�����ot!��r��0�\�:LR�u��lT�Y���A��'�.he��c[��n�⠻��Q�|�.6.��Ou;�TH��L��6B��r�׷Mr��B,`���#ju�4B�@!��4Ha��\��N�&q��\"��K@Ό삌/�d��Bc��}j\:;H'��U��x'?��������E}�H�I�	+�
�}h�M�&�e"Ϸ0�e9#g��%�!��)\/��n
�}T9bw���y،N Z3�5zqM^���n�j�6���� +��XNG����b��;��T@�a G�*ȴy�3�R��ڧ������b�S��28�b�x\�'�u�]� ���� ���b�1mU�zT�R��ds��(a�A[�	,�X���@�$�7�Aj|H�_���U��{��S"{�	�q�|��+A��C&��1�&���z9!�K+�IןGEg>�d��u� �%�v~`���Jge�i`o:�s ##�o�&C̦��M�+�o��1��	�ǕyE�U[�@Un�&N��%me�CKt�) ��b*�X [ D~�G�o�����G�=��G��z��l����<.�q�3kd������MO��~o?��w(�Ckٱ�>Q/n�j�aإ?\5�P?h?s�[�������Q7���Jt��b({Z�*��t�a)e��O�}�f%���JKe)ḽ"oz
����=�A({�3�k���#���2�-�ulߘ%��v�U�?��Bg�8N���_��<.�3~\5H�AÉ���b=[U�ҸO�F�'���`5Ŷy���(<	5�c�u�?pA$�:A/G~8��:������@��d�]Say<ʍ�#��Œi��K�X��~̔�����y
��� ���x�p����~&D�}��~�{� ��=�[�?�,nt�U��7�eWT�����ۯ�|���:	ǰ'-�oA�g�G��aۖܶ�e�¼$pr��KP�S
+#O9�*���i��W�~��Ո��F�=��dV<nb��+0�������F;�
~�X�lyZU	�n�!F��}�q���R�HѨG�iFc0�I�������1!H�7N�R����� �P��zo���b���e�G�LS��|���*��B�Z˸�v��e��}�2���3S^1��r����%l�L��/V5[��64�����l�B����\M���};@ć��,O���֗8-��/ʣ��z������P%Hx~k��c�\��i�e.X�$�s%�A��a^�AE�=V.��N�'H�R�(W���ɗ��Ԗ{��-LE��bLER0���N�aܖ�Q������3k��J�)�%�fHr��5��=����,����d��b�2�u|��%�����J��`��R����3��4�C[=쭾��G5g��cQ��b�}�m� �9uҶ����H��5 �X c:��w��A�-0O4P�^w:y���9�
^��@T�i}��ѧ�W�N�UnL�0�U�֋ǰ�P�ر�cչ�?��p��΃��n
Zm)\C	����F}0�[a���iŲ3$Ct��Ԗ�L��v2n������\7:_b��c��A���Uv�k�9V��zЁh��t�A;��F�'_h���؍�H�D�PsY��9ݬ�53<�y7e^y�ù�6��d�׏�W߈E�;ܐ�o��AbҤ
3r.&8:۰|����������>�t�]�u�@�p +���vW�f��#�&QF+����׆�8X.#2n��ڞ���N�as";����Y<K�Ԗ�TV��i�J���1����� D>�C����>���h����k��}~Q����(�s�pFfўBh��7�&��U�0�]�)
_m�vr��fd\kI�_S:CƇ3C���?�&�2���x��?��L��HNp@Qh��=d&W' C���(��tjցAlP(�r�,�
�����g�7�`r���΅����&R��j��
6�]p�g�2��77�G ��b�}��nꭸY���{�?'XHLM_Z���_⊇0�*H�m��c��R�ww BQ�.vّp�R4�T�}���x8�*<j�i%~$+I�ئ8yŎw:� sۂŸM��]\� �Tu�o���Dծ�>[3=i?S�a�涭	O��q@�����_`��گ�5�<֌�o*��˱?Z�[�[1�x�](?�q���5No8�Pgk�m���o����6��
3�g�Z[�W���vŗ`Ƿ��BcI�g6�!|�Q�j؀Çz��l4Ȁ�����;_��݊�6]4CT=�/�����1���?@�\�8@��/���A�P.Ϡ�yo�6]�*�O0�Y�K��ۙ��9�c��g�\�A��hq;�?f�d{Ij���n(�w�<<��c�W��̅�MO �/	���@�g`Z�a0^:Q�&m۵.Nݗv[s�mj͟,Bf�|�lJ�jh^ b���|)/�OmS��^Eǲ�ׅ�aR����7�t�� #�Zd���X`��e �b
��m�7'A���RF�K��U�{m3�x�E�&e<���,E�k�����)+'��G���3a�(�F5g'�iBʷ��]�����."��/�[yd�qE��%��=)�4�R���Dr�܌��o�����*IL@j�ƕ�;+�Hf�/�4c���zAo[�=�{a9��1�Y����N��x{�zE�A��^�p|����^y38+��-RZ�ߩ�C�2>�,���M� g_��@��3��4Y�����)C��j4��t0���_����"M:m޳o��oT6�щ���8��篠#��<�`y�BkF��-X�Zv�%�Nq��ӛ |�����g�ׅ�G���\�:O�1E�pN$/`z]���Ǎ0�g��D���)5=�Pp��N#�W-�'������-��t�
d��)�U�"-��0"�>�h�$�|�xb��>���،C�rR_�B�;�����=�4�4�}�v��D�,�`��R��gե��f��W��"��Q�
�ФQ"8��OQ�2E���җ:"@� R_�+�I-�)7ꭽ�C�|��fB@P�tOJ���/p�9�.B����ԩ&�E����u��D H���L"-�����+?�����N�'�rm���0��ͤ��0ؒi�A�I��Ӌ����/jD���ac�z�?�Ʈ#�r��;+�8��`�X;d���R��x$[I!��שe���F�+�H�R�	���Y�c]\��C�i@d{�3�q|�G�������q�,<�Q��}��c�U���j����|b)`Xqi��Y�f���ؘ�j�+6��䦾���KM3��S6�#���GQ��J��w����M�T]���@��G�����a���BW��Ʒ�>�`Ƚт�f��*�P�u�zi�r Jϭ�i�ϝ�~P��m6EƁI�Q����4ث{Z5UV)e�qҌ���3�!ǟ�A�o��!hi���y22y�r��R��~X���̤u53��ȣ�@6W�\�-5
N���F��*/�D�ȯ��?kb��� �$�5Y�݅D�-���d�`qڮ�9�
+�1A����8�1���������9�J�D�x���`�����<89%�1�ɟ�M��@+�OK��u�LM���,���92�ED�S���mX�h��9:v(��dS����=}�p�x�4�^:x�u��RV�bM���G��ڝ���|�|?�#F:f�g�Ӗ�2		P�<�?���7�U�F
��?�+�b6su�zM@w��k7?}]�������4A����[�c�;�ۡ�B��IUeW�킰��s���ۍ�����ae[8���FY���Cte+&�;w�u�o�� �_�]��h��AՐ#��WT6�X�.�b"�n�TΩݛ-uSq�T.׊\,��W�+D�}(4&���Ƿx)o� �~�i��@��-��p����թk	\]>Ω�2�d81{��,s������[���K[*umx����	����!��~x__����XfɌ��K�x�C��o�eE��w�B&� �h2�|��Fc���L�t�q�=�b,Ql�t+K���
0F*�2�/fm�(zs3c��~��<�Lu�Y�q>�FS�ȑ��6n�̹�~}�.�d�� nٺ�|��rt߮��[���ՄR)/��W��s��x9&�)��Jm��[�Rs���+!W��)6�(��[��1z_�@�kMZ�]c������A�m�cܺ�A�oL�NKr9 ��BޏF��> ��./������=7�8�B�����ѧS8I٭���7�6��g�Y�12���5�V���+��C�
�`� |*�}<�^��b�@�������OIy��edA�b틷��j�(�p:d���\tp5��D�B7Z��H؋��Y)�W'P�xu��*J�&2'OQ�q�\D�t���������Z��H���D"a��K?���E]���4���p8>�M��}5�"��E��~���%�J	�Է�H��G�k���foewU�ħf�z�jz���nй%nUj?�w��z$�c�W���jR%�wTԻ�M����E�+om��7Ƞ�}`�7���^\�9�s�%O�q2���y�{%��UC3s���C��"�P\=�3�3S�����S^���<		�7Y�C
D@���&��Q�(�9��W�h"�E =���?�L�vbP2�#���as(m�3�¨�s��4��z�;+X�E�lO�[S��X���h����c��w!�}}g����Y7U���҂>�Wm��������^@�ɠ��+��:��]�l���6��P+M�n�x􄒽VkV/��\��X��(�c�J3%��~R{�|?����fI�$ۛ$C��2%9���M���O��.�?��Pi�*kB@���v%�z�DL>���D��!��х�#���6��W�y���4l�������l7���0Q�4MyCkJ�g�d� ��O�Й�����ʉ��"qM�����%�r��f�&�ꂌd�kd�N���$#�+Q7�}�o�| 00?���P�?��[w�*�(�Z���χ'|xE�������S����T���:��q�dYW�����q��G?� ��DM*����n���+�[�1 J\M�Fm�֜E*���3�FY�M!sT�V�e/]<��JvH'���<�!.���!p��j�ǧA���<!}�Έz��x,~�g�qfVo��WD���$��4�Z�0����R��B�~�.�@�o�I>��`ո�1�+�^��P����j�^�����2��Krt�љֺ��Л��L��O�'�I��b��kթ}!�� ��p5���t���**�y�i�F��s?2Vj\��<�^�w������󲵧Ӣ(P��%�[����a�e%zX	"N�\VNs8�̧߃cA��mȚ�O!2=�̎�'���h��$L�X���4x�������k��'9Qw�1�.^n� �$(=+���w՗�I0�Xgnq��T:T������s����#OPS?vZ�rO\:�D��x���/��,�N:t��a���6Y����5#&&�_?&<s���װ�6Y�
�q=5&'vFff�-�/��6
ʥ�����
���tM!MKI9���(��j��K�]���@�Y���>��Y1ps�K�d���ό���Q�E���B�_���H]�G�+�77&���oU^.��U��Rז��ۀG��C�[�r7n�֠��;�+d�
ht��4��6���J���F\�K�9G�lN����V���5��]j�%1���ɛ�.���"�ۢ:�/v)���vV̏{��is$��!dP-��O�+��ќ�-$S:�{9ULf��� �\�ʟ�0��f�����/�c�~J�+��U��㟥�|��s3�v�9}|4�ϣ�f�d<33�ڿ3t@d����8� )&щ��s��{��4[�Pu��Er����ױ���� }�94+,C��Y�	����Ӝ9������RnM���o�U{�k9s3�T!��Q�|pP��,���LO�'�g�sf�>���3\oqvw����|C�%*��*��!�;���{`Z ��wj�����.�)1ͳG����k�����
��Y��B�����r�4��[x�tA�p�9����Ȍ7^��hmVt�ciT�;"9��e��h�ad�_�v��| O�)�2���3m֘ %59�Ec��sC�����(�[1 �L�e�Ő��5����NF��o֩����]r�{������2���>B
'����8yf�y.�� ��8���Au��)gTc6i�iMLd��s-g��nPH�}����މTs����/�1䘧R���Ӌ����4����ԍ̟E��?�8K)HY�~�a/��c���P�Hy]]VЄ�H�N���rjow��XP�"�Ͻ�&F����۟->� �}6 �pc�(�3
�&�d�"��u<��j` �E�&� �dv��v�{�j{Y^n�K�2��d�����eW"ځ�IIE�,�?��v>�|@iܟ��h4��E�]�w��Մ�T�KF�a3"]8�>w�"�t�A�I����`&R�4�G��D�S2j�^-V`wl �wi��F�!��Q��Z?�F r_�l�J|
��\�\�D���
t
�Rhp�٧���k���z��[�v�W�A�FSe������	�{ƣ�I��6"��<a?��zR9���Qz��*��%ԆF#9u�^�h0[�(�et�]Il����<7�6��8\�(�ҟ2����^j�>~����,���J���)�`I�M[@���2��u������\Kց���c�Mvv�2S&���2���l����9���t���n��c*c$����-$�,�#P��AڒCc�r(a�g��V̱G�U�k)��l�>�DW��!���{xqɤ�3a�/�ɰ	6L��D>ENB�rOV����ب�JD
ǁ�w����Zۼoޒmۯ1�Vw��Mcz��%�1�PX\E2s��4i��9��c�P�� k�Ȃ��z�!�*�����o0wo����\Рh�O��V��ƀ�
R�d*���;����>� ]��!�ݛ�.�j��;�~a�_8����NY\O���I �[s�B���D���(G��PsJ�51��o��ޟ+�>&�B����5{��;��%�͜�̕6>�2 ���R�o*In����K\��M�w����
��m�8�|��-�wT �:b��q�}.\���4��Y׍+H�����ȴ"��q[�ޜ$P{��P�նx?�el\]gV7�ҋ/�\���͜��[��C�:HʓY��k��N-�	#��zQ��U�|r���؆���E�7�X�Y ����JT�>�+�D����F�U0ϭ��N�H���R�Ob��#n+�΁����}Κ5�pHo����~bp�q���S�`9�l2՞.�A������Y�ν�,b��9j�<��S:�4Zs@~v����)�KG�N�:�=sU,�a������oh�A��~}�2ȣ���7�xbL���.�6�G��B���~�@E�O$Z�M;��#D]�Q��U�+iMC4�K:�2\Å�TA��2vp���v���(�U���v���g6��'�!�Q0�Vk�y�ܺ��<�;�'M��3?���JG�)ت�k�����a`��p6�;�I�$� ꩚D�$�U��� ��8�'�^��D�)��X�8'�ߋ?�x��z�57�����&mD{R�q�r�"��|O�*]g�Y9�����$ Ӑ�N�1@0����ض���y�>��f��q㍏�G�6�Z�Ns�?cS�S�EHIpϲ��y��W�Q�*���sѵ��
�R���м�g�/��	�8���_�^"���r o�b*z�dƺ���u4�bJ< �qw��wY�]{�F���u� �iՃD���)��y��kv�h���L���ާ���n��e�+"�[�a����a���8��B�+:�b�C_���.S:��N(��ռ˞�z��������^�r!c�ٿq���1y�D�X�-d|$�5�j���`���8�t��2D�;`��asr?�@�U�B���}��܊:`@Қ�f��\�tL��^��3�̳�e|��%z��Y�OXe隉rԚt����Ԗ�XY|����븤�Aѭ���T�$�g~�D�R��|+u!䶖�QD`�$P�2���-?��"���JV���#��"�� �2`�2��Z:T��Ǡh-���xYF����u#}��3�e�>�C�֋\��;��K��ΐϜ ��q�&����+�&���bSl� I��n�(��^��C5Ê�O2 X2����3��l�m%T��Ξ��~����ũ����PN��VF+p�DOZ�&+M\-��2%�}�Э)Y/y���h��,��,�R�]p��>/f�^Fk?zt]����h�1)�!�i�J��Sd9jS��&\�a\L�ueG��2�(�����t�b3�=6m�+з:����փ�̍3j�}�v��7E]+����{�\���<���\����}WN�&�U1����� 
}`�ꊶ(��'b]a���O�$�]�W�sy��J�:��* !�H�2��O�]�v�{���FR�˼�m���4�@q��N�~N��c��#��~,`���uϐ��b\`����!��VxT?����X����B\���|�$#Z7f�m�XAg��@Ղ����e� ����;h~2)��%0 3�������6x���C��ɸ�JvL:�;�!U�����u��kص����h�[����`S��1��|��!��rC
h!���bHcg{���|sTĭ� /p5���)�#�DjV)d$�ܰ���0_��֩�a"����'��t�3�yL�cح ?+b=�Z��d�g�$Ö�9��}Z�t��?��� ��<e��B�ɼG`ր(ۋ��2Pa~ߟ��`�}��p�p�ZV��� �G���aMį�5$��d��OQ�[Q�K��Q�a�=�(�����AB?�;�5�P�
Kq�E��BUl��$�v:�̈́�V௄P(*�惪r��w��JA��aa�������=��	:d�W��.e��ĝ�>}�o$M��W�. ����r#md �`�=��Oڪ��
h2Ӑ�䬎����1�1vr����H�� Ѓ�b����N���]��O%8Ӕ�Ś�f��R@r���[��3��
<��F{���n	t.\|��O����3�u5j[⠽y��~��%���3�b��N����)׻�o���C4~-��b�C�0����k�]7���"�*
b�e6�5@���zx"��⎡��h�=�/���T��Q�N5�-�Wߺ�&�8/�5D�W|�4`�W6�q�=�����ѣȏ���/��]��4���j��a�
y�~���4��$~�(pa�Dr�
�5>lͩM�y0^�I�����R�/�ۋ�7�'�V!�#"��"E�{=Bhcv�3�KؚM��g�zn�[���n%x��N��ӳr6�=8:�5e&�ws)�D[�g�=%C#��:,���V;tIbO�7B<%�ޟ,㮣����'��A웟z� B;��>�k/�kW��._ss�v[�v:r �NV�9�Ж �E>g���#x���$^: ��K}`�cX5s�t!����di	��3!d�e
Dt򊇤v-Flo��Gj����@4�l����L[l�@�\L���lq�|ASȎuE�hN-4$��-<�3�Xܜq�j��f�eH�fttE��C�p��V���"1j���#O������&���<�Y_�ja��M���R�s�cR��ۻ���V|��v6�q�lt�j �̉��1U ͝h"�w��\Ui;�X�����$��,�'���jt��FYN1N:0TO�O���c�a������I��4��A!�.:�˾Q�RW����6�� �|�E����skCT�7��bܟ�ZH��c�������X��%�޻���x5}�C�u�yii�I��x���Ǩ)��S� ���+�#6�x��ه���2Zg�񪝺_�C}M�8�����v_��
;&��Iq��1�Z؟ʵ͵�j����O���z~ڳ��4�bޖ���Y�a�S�����I�,)jف�u�2�A��4��׼�1^2mֈ��1�s�E��������q��9�?�7P.�#�BvK��r�N�s��<����;�� ஓ��'t�l����L���	mn����*#O-S��(����]v�!��nU\�U,#�������'t�Z0H2|]Ϋ�'V�G�W�V����p+=t�0�-�C�3���
�#��Z����H�v3��Ű�|(]��f����C_�=�}�^�7"���i6�����Q�fB�
�*���+;�TDy�r杈�c�${��J�� ��r�p�\�]i����t�W�y>cڒ�U'd���y��6�c�*~�x�=�a�DS����Ѳ�a�Ҳ���-�=���� ��sX>���sڤ���q����N>������m�N	ޟ,��#��(7��10����]��+������,������̊⺟z����Պk�/VǴ�B}@=�_*͂ ��;�������?�q{2>en'�-A�7p����z+��IWo	��-�nN�j(a�ɨ��a|����ST����:�����-9V��i���g�0�n?�oq�u���f���ʅ�z�?P��p_D���hfw�C{ݔ��X��\� X�ʨtx��$�ԑS������"���r�C�gd��`�/=
�l
yo�Ϧ��t�Vj�?S���,7�v�/��K<i�{N��!FS����N���,i�S�S��k5-qG9���0#"�Σ�Ga��tQ]���0�knп�]@ޑ	|+l;`q�n��3��`2k�^2d��	���Jf.!�j��,?^�p�WBn�0��ot��MȘ`��N��{�i���vcA7�V�A]�7�Tx����Ư,�;��Q
��>g��9�Z��í��4��*ٜ ����h�
ޕ,���`�wS�ƛo����f���\��6f\=�{�v_s�WԄږ��=�`f���b2��U�Jt�(��(*�nJ��5I�LS��l{偰���Z��@��"��\8�\d��x��Ǧ<�6��fw�~�C�:�K�4,�5�1�4�JE������t�`���Y�i���8�ΪS?����,%`�=���퇕/�o�X5m#!��=�����Í^I���,�'�n�8: ��|#1Lc��1l��c�]K��y;ؑ5��V���VI�d��}<
�!&�ی�[�"�p��|�흻]ձ�����c�J�Xc�WM�xY�4�h8�
HXjٖ������Ș���*� �c����Qw�5��W��|B���������Oh>����*����+��B[�O6�f�����c p&_�~�i"�A ����T�W��yo��Ī��%�!���~���M���u�4�]У���@��� ,�6�u����ks�Yf�/��XPIT0XM�]�вX��F�1���	����J����G�X��;����͐s���g�]�y�aO4�1
���n�Ub�b�`S����PmU^��Ǚs�L7x�m4K��@w��c6۴ԭ�G�3���䦰�*w��
��9�c�I#'�Z��H�hd]��蚊�^�I)�]:d�ECf��ȴ���hړ�.��}ua�\����1� �hG�v��-N��3���?pk�ĲKY����]D��*)1��O�7���)i9�7J�	n(DE<�J{ĭ�o.�;CV��j�`��v��I��_JZ�Y�>�H������뵀�W�8��^{7
��QW����>rop�h��Z)������0@��%LCt� ����x�����l��Lo�SA��z&��Z���k�;�v:}З�#�X�j���J�L+|5jM����aP�㌃l���*D��.H���=�b��
���:<s���"��Cߕ;���+j�heZ�LD�1�H���
`�.r}���Y*��I�ܧ�ѠKe�踊�`w��l���|_3�5�p��܊)K�"���8�*:b��p�	��ŕ;Q}��S�p�Wfa٨�J)U���4CB�d��U5C*�j�W�=׾�V��/�F�Em��@f��W�)e�e�yf�G؈�\�!m
v���'��2SD$4����dm��n�c'D��6)N������u:�:մ��*Lo�O�h[Ͷ7.���U��OS^���1Ű��j��ํ�!�Z�GO;��z�����
!X�V� �ٶb��˺������i/D�Oɴ}�Fib�͞)��> rh�1g�/�1F�lP�����	l�1����L�T���`%��~���b��__5;2�G1�D�u��1�����7���CM�sg�_�h@��w�s]Ki�83~�t5�)�oc@	,��h[�?�'t�%��i�v����Z�v�}��:�]�fys�%��\��͜�j�2P�wG�]�CJ�fV����^�:�j��H��]�����	K���+p,ba�zHr��b�3�w�P7)� ��V�t�cZ5by����851���Q�ȝZc7��
 �4��}Q��g�mkcbV2�"���5,lՔ���&�҉�^PG��<i#>C��[3���؋q2� &s�����ƙ�F�H�*�5I���"��2��5n|�>���j���uرUOI��9�����nte����B̆���������*p��̧k(�����G���Q�|hǯ=���f�2�~S�*O�w������H�m��H��5 4PI��5���£,����:�@��VP�i����%�P���B*`W��<`7����S�i�f!�i�,��a|K}�}M���3�.Բ#���R��ȩn�%�;�M�Ȑy�|GK��r��iՄ�O�I����ǰ�K�A���2���}��[�~9�Y���Ѧ.x���:KI�Z"9Gܿ6���4ו�a0aԝ`+�N.��r0�WRĄnG }���$���)@�����T�L4�`�:3�'���'��At���t�Az�H=�:��K�����$�.Z3g�&u�u)���'�r:Z�*�>0:SQTG��]�٫���u��B={�� �$w�_���XB��^�7���GM�!�`�E�6�[�[6���.��m>H��X�*�������c1D�,�� J�>�R�B5f�����X'~�ȋ�[y�ztpӝ������B6C��[�Q���$!���o��u���B�GZ��0�hOi�*%Oỿ���93�ߤ���.U�W�$-�����LjWk �N��K.��D/;TI�m=W����<0� w$JhU����Ǩ�g,&H�e��Õ3��q��Y%�_�2�՚��E�+;��D����+�^��e9~� �Obd9!;^�Q�	�4���)!2Y��V`��4n�``��8n�d
��Q2���v�!h�T&/�s'2a�0�Ĕ�w@=�H�����rv=�D�H�)�~_p�����{��@�L��=�L u�,.>�G۔��wd�'H��9i�<0�CKgKL��#&O8���0�z]���{sw#ō)_P���)�a[��P��fs�*moM��2#�@��C�@��g�KsG8��V�Ij��J�ڭ�jM�	.�Zb���x���_��F�"h�����#���N=$
��F˲m;�7��3&���/U�m��^�@�-��bA?"$	�������]���@�C�GӒ�Qn�'���/����{�@�Nj��2��"��E2ׂ� ��r�Ｋ���[;<_���~����T&Ą�G+�v;㻨�);��1dV��a�f	�Ѝ����@.A�D�hP2�x�zHcQ>U���C��W��dNj�xd�Z<ޓ�$C+J�Hi�:X�A�?T��GH�����/�eXʝ�����C��oM��+� d����~��*��Z���t��)L��0̦%�	;��b����%�-*#r�����6T}d��Űw�V������ؙM1��� o�}��M��F����W�CG����{������N�m}8ؑ� 	"R�'8�7Ɛό_-��GT�=��Fl��M�UEЌ>15f�����A"�Ȑ�cU��[���N�S�sXh����:�������߀
t��!O�v�v�@�U8�Ud��.	�?�9��B[�[�d�k�P�!7;�"s����x�8\����5��|�cf(	b��HY�À�d|z� {�8f�S�����U�#T�w��p����0|;��װ�t�iӿ��v�ab��ڇ���|m�9��>aDC+��W�3�bn���%��|��WW�Kv�u��p�q"�J;uF�5hD��\�Â���Tfa�[��^��ܖE�WMԬ~@ǹ�仫�FwT{Oo���ge��ʐi`A�bx�]��I�H���>�M_<��$|s���Wa�����{�I��X-����+R��N���I���Ⱦ�+Sԏ���PQ!�W�%�6Q՝vލX?�4(�ß��V��kMw�A&Fr�i7�R���@��������t�_�&:�_#04�^'�%rn�^g(�\����Ȱ��3�*�G���ց��1������j�4[?CbL=�D��L��s�3<z�\���}w��LS>6l�6���.��G !������`Q;t>�h��}�]�<:�(8c>�G�E�ȋ����-)�P��1�����J4��y	%O�#ŭ�����n֭?3�:1�5
k�ኅ�\j�5���V�g�^�3�Z5�n%��D#��,C�I��#��t��xڨge�����5�b��{oy=��2/ n/Q�<j����a�|E4����^�F*MQb�����ō�Ig��˷�R|D!���Ҭ����ߖ(���0�sEf�|qq�R� �\jv��t)5�E��Y��8`HX��F�ǮUIy܎���(�:���7 �3�C��DF��!:�H=��]�W�?�!��Ւr��I N7�×_�_��&G%���fplB�w�n������X3�oX�������ƕӂ4��.����?b��J��*��^(z�ee�kH����(2��މ`<��@��B�����*��bJU�1�-V�)Ǫ{V 5��w#��s}X�!�-ʥ�1��KK�P�� ��LkWZ�h��𚼵����s���P&;G�l�Q�F4���,���<�2�����UZ�oֹv}��<˯i��u�/����E)�k_��a>yzO|��
2�Z�
}gT4������i�Y�pj4T�5��&|Ӵ�1�iN�Gπ*�8(dzl1��$����9�V��۴ƴ�H.3��܎��76 �Ė"8��{Uһ��A�՗pd�0A�������ŭ���2��q*�����M���ΰ3��
os�l/-�.���p�/w*]j1����� �Va8�l�o9j�u��LjٖG��ǟ�W�W���lؑt�#�@�X�}b����\�,�ʿ)��
u����$ʚ�pUs�����>{�k"�9�B;�	@P��I=չ���B�`�Xf�j�O~��5V�W����8�P:ω�K��9��� �Se�6�oV� +�w��0p^Y��u��?�J<����ծn�<��(�t#T�k�k�"1ѿ���T� �̷�{�44���f���3 ����s�E�IO�Q��*D@\���-Y����� :�q^�c_E�B�U��A�d��kǣV�*�e�"`� /�u���Od�{	��f,>X�o�c��{�Ohx��;p�ѩ���7�'h4V*ա�3{�s��_�$�Q?�,R��Pd3f����j��nd8J�����DX�%���P���Ix���/�-��W�/x�
��޽l�(�t8:4Z�:H	���(�
�?��A����wL��+*/���ϑ�Ds&�v�m�(4����������Z7FmB.��U�0����PqBD���V54#	3�r�/���o$3��2��`�`*�ZvT{�_l���gX<�<tU���~1�z4Z���Q�*mM8�����{V3�:J�h����U���m����z�I)�y[�5@?'�$�� �Ć�����6%��bK��qDҞM����G�����*�{]it�u�x)�9�^�Z2�c�9�(��7m�n��`[�28��w~�l�P�|j�.w��[�A/���X���$by�T\�%jB�&t�]j���<.z�:�#�gΝ���%���>��&��<X �5-7�F��{��IB����\A�q��@o$�3:mr���#<לxQK=�X~Z! ڎ�^$�f�hޮ�@�&L0	�Z�?�NW��7J�"z�c�� � ������6�U�����p���oj�k0:�{���gnb�Z���+OR�o�� v���h�L�] �af��;���s��Z!�v/�ַӦg��������M#����xKG���<ƭ�#�;k�EFGbj?�X���_�SW�^��ťu�J��=5P�*� ������b
@�Șif"D��dBn�����e7嬪�X\a���i�0@�_��\��ӦB���n7~�*+WɁ�:$d�ri�G����Vŵ�A����Q�2�4�tp�ܲ��a8}�Hp��]�3SښvMҠ�M��i��ۆ�n��O8p�8�tl����
0��#��籽RU�מ�d���3,XT�����g����w�߂k��>�&��2	i."z?n�EP�B]��A�� ����7c�pjě��4=d�e�g�ƾA�+�񑜟��j�����;����7K�AW�3��u�7H�s볝�.��_ʓ��T	�9a�U-ߪ?�yN��X�K�k���ϡJq�DPϷJ6��f �!Y��K�>er'jU���jt��gn�In�'��qЛ�W�X�nu�b*������v��-֬����A#*�� U�[ǅ8����p�T�n@�O����A��_ ������zU�3����-p.�c�6��,�F?�[T؏��E,a^�)���3����$ؚ�*�?I.�4�A�<g�z�����y��&����{vD�x�b�[qU�6��_�%%#4�Ӽ���<��Z���W���-��8��J�V���n����_�8R�L+6�W�]�v 9��S�q~ݞDϸ_�f����T�� J��~�s!�$��(=28��3Q�8�3�:N)��@T����F���)x�t�E�_i�j����ܳk��0���ĮY/S��S�؁H|�Kir�lf�A5T�懮g�NZ�&�k4qH��������>��v��r��T�;l���v��w%|��RU�w��P�^bi��g��|�]���sB��B�|O�O$`�mnZ� z�a��̞vǬu�����+W��D���6����4?\[	�b7��}���X� bF�z3�!�v���;�>��� �D*6$u�D��(Y��~���7��LW�����o ��	O���Ø�s�ͨ�xP���p�\��c�У5xK��=�M�S�gҢ2���Z�S�Sܗ���MK·��ml+d2TZ��M��s�қDM��[ky�gٿ�$MlM#=|ykX�Y�>�Q" ������3q^.� �Q�뭫J�^�d��M �;��$B��=�Ohxj���r9 �0W.�:3K�G��7=��5��� ����!��X��uʼ��[�ʯE$Io8=×c+��uߟ�`�}� �� &],s�����j�\é���J#"������8uH�y��U{� a)F~T�+�>2k&kHrf%4�%�U��ʹ��je��to0���6�nz�wA!߽���#mt2�"	�r9��g�:�9����>�Y1��X(���8]�y����ųڇ�����fa}�#S�a�d���['���z��*��fT�l��W|1H��aW"���k�I���-X�wy5�JE�N���N��z'GY��KM�B�涜5�����2�����؎���N#^ ˲����f�a�h�R��6ͤ�]Bn˔ʵ�􅲲�;�[I�t{�v���W��\�"���]g�½�[���r�Nwj��:��p���3rx��;kpwG�ۤ>�1މ���	���	R�d�ؗ
�-�����S�F���m�fr��^�7�G3�c�ofU��_���b�Ӣ�}����Y�d���]�my���vcqMa������d谖W�l�+b��(�O
Z��l_e�}+�n.���S��]�R5�&�s��g�}CX���h!��%:���
�����"�K]a^��G��e�Z�6���-v��iY9̠� ���~.V��X�4lr/h����O������7A����M�1Ǒ�U�	Pm#n2í���'4 ��/���'<�\��_,H"!����xJZy�޷���S����Xxݏ�:�(�5X0.�O7���"Yv��q����._೦r�Du5蜍����u;ގ�Mh�z��B��$�ъ�tg�܇9/_�I4�Aa%D�(8�>;�6��
�@q[56��*�f��IJ'T�)E_ժ���U�� ���Ӣ6u��	��s��ϤEO���я�?�4e�߁�n0/��fFgW�.7?��ڥ8{<�&M|�1F��Y���u��$��J'tg�Xx�|�]�D�z1rAo�Z�?=D@�O:E�z��r+����Z�zKfa\�1d<�T1�5�z`Es`�K"8�w���I�5`� �Af�MSOy���A��t�(�s�ώ,�P� L�ٵ�(ء�
��=K���fioB��q��v�d�:Eѡz�8����(;�=}I;4��� y������c	�X)GJ������ �j�-������@��ܘ�	�*��b�/�Γ�K1s��E1�{жW��u�
���C��Mw�Ae�x�,����n�k
�s��"f�O��ֻ�h`̈́��j�w�����j���N��PV�p��_�y�	X���RJq� �bE�����O�.�E.�N�X���9���v@o���>d@qN#+�/���O�<�����H�^�Ni������nD��Q�bS�N�M���E Į����T�}U�A��g>5�jaN<[I\<��7W_0�S�>��� �G-OM r$���wҔV��/���2r�K#z��;�Z@Th�m3�-VA������ ��w�
�>�=�ly@�3��,'&t*��l��5�j��2��Q(^��v��֪�sP&5��ok	��+N�*��"�6��m*SN	2�BE�p���{�j������X�(�Ĕ-�����h\�X��$.B��-Z0�z��'�80�Cנ�_�*	��R�5�R5�� �����t�u9�*Z]�o�����hj���4a�o�ѮVמ��$RQfS`;1�.O�>Y��+F�I`	r��~��Z����*&J�+E�W~Hۻչj��p7��Յ%��Ekr����<C����ѥ+Iu�J���j��.H��yZ{,.?S����,}G����l].!�M�Ha�n�	a7m�K=ʺ�w_2��������vg^�%b4��J�#=��d��KWĄ6�L���ո�5�d�u�Vč�Δ:tN�]7AI.�kYq�J�Z��]sH�L��zb�:�0 ;��Sz��B�/!��$�i��i�fH�>��O����ӥ(�����t�TQ83e�<�� ���ܗ�~���0T$�C��5�\Y/J��g!z��GR%��o��"Ƿ�`o�JH�bc�9��b�:~���I/��<��L}J/�Sa�i��s�\��n���a�h�:��k�s_�� ��+����7������~��\�X��֟l(O���a�V&�p!���`�X�=m|��8t�����<D�I�=��g݃����|��~�(�?�?V3;��%Ϊ���Ĝ��s�o�w��o�.�-9��8����_g��X�a |Q�<H$��� ��e�N�;�c�؞� �7���P�6�躐o�@ݳ�!Ao�����v����v/Gv�n熩Tc��/�.���~M�S��^���ʷ��|��� ��_Z��)j�g�-�%�ˁ�ul��w[0��@1�|�qhc:A4S�|`�����?G	Y�'#x�!S��ZW������c�V�Yܿb�Rf���]�_��}����;��$��TY�6.+��m*0��<���� �Ot2���u�B�؛���!{�l8t.�6�%�M���<���@^�d��H��QFչH	��㳼��%z�����?�s���9������ �:Z��y8���U���	v*yQ�ͻ��
v���ޢ����c�vM)5DL�6��C��\�
[)�H����D\4�Ϩ=�@F�n�'#���u,D�MfP��]�mx�pW�4�o���)љ��Dh��OrO;�BYN[˘ei}��^[YT�=���d�Y����qUe WT̢�5{�|g$��-�O��ZH)#�.YI;��X�w�5k���S*g���8v¯�n�Ձ�л����kR�h74JE��i��MT��0�򆃩���'�w�X�z�+q� O�󉝅�����4�Z�>��@���F�V�YŔuֲ*���6T��h ��yǈQ{����3A�'��;)���뉶K� ��)ո|��ZO�Y���^6��ѹ�I��q�x+��D>���Pdu�t��f�j,Ǻ,n��.ADnI9�����6�sb���L q��~BY������c��e�\U2�[�rRW�6�{��;NL�a歴����{.���dA��`q ��Ob����Bևc�"¨*m�,���t؊o~�$6�5��cvQ*ɭ�w3�%&�ʸC�U��Rq����S�<�s�o�����W@&@�o!�F�2�7CH �՟���)�h{�['z!0�Z�|��)�sq�o����f������=���� "Y��^G���_������t'��|)Z3��5���E�E��$챦Fv`j+��qZ��-a�
,+N��H�I�[��B�n�WV�����1}���G��5��\_�!�mI�X��wD�]`��,`j���`ing��p'^S�	^a0�$.�$�e��w�7��L&����h�Y�R1�yY^�vI�R�߻�I�	��1����c��i��`)��W&ӊ��y8��4?�K��'Go�3�� e�xhϟ��'�3x����[�$q5���\J=]��%,7�/������Π^B$��XO��[+Cnq8�8/�2�V�n�?�T sͩ���ʣ����f�r%�(��$�����g⅖���p�t$y�Om��&ٍV�+��k���Q畹!��ӽ�ى��]�%R��G� ,pVIQι��(oƊ�D��)7v����恺@o\�0�Qü�e�Z���s �|�-d�*����a��
>�˧�AK��g�	���hs�(�&K2�y�w�V	��Fn2wI�ߑ.�S�{u���3�&����N�!�^V�54��7#��F�P/�N� 5�C�C���e�p���rV1��ޅ�+j
l�iy���+p|���И��i��6�2=F?#uG}p6ec��`��e��<ȗzI虜xo\�bKꪘ�� ����!���ׂ�T'R5(@-��Z�쎖��k�f��J�XȀg���n�<�o�RA�hԑ"�k*�����07����~�𼜍�O7)`["��zי���ⱴ6X�Ծ�c�����E�o(�7�4���S�Ԑz0N��e��٦� ���Q�y���XՓ�z��c_��{<%f����uI��&�4�X`�{���������P(�P3A�q��Q9/����*����������ړ1I<���'K��p�O~�h$�i�-�4����O��Ð@�A���$U����mH�����@�E�>�6���e�����K��o�F�2Zm"s50�~������^��lo|�)b�L'�N����}�Ǹ_��� BR�G������]\i-Y�u��:��=����HJ-�O�x%u�$�G�[�2�)X �+�f�8>�G��.�B,��|3���CpQL[������d�L�q��j+�[��kat�Uי+�@���y�d�V�<��J��Q�����@�q���i����� �<y��f�O���9�(��5�r<M5�j���ᄯ�F�>��	�r"Z����nb�k;�ÑP���ow��W�_(8'���)|�1Tաw�������%�c�%8L�L� (�.i��S��^OiJ� �=��R�̡p��B����k�;��g�g}�	�H�5�L	at��5��c�g\�,jT�ȍ����(c�UV�R���p���io�3��#��"�j²�'ʕ)��>b�@�܉�'� ӣJ^�����MBo�Ʊ�� �x���B~�cl3�dj|#�l���G�P��$Aѱ����m��q�r��`�k���15��<���*h[z�H�4�{�O[������*dRH�6ſ�S�qhX�#��WgՓ����p�"�%��3�B��!���&
���Y�,q@$�H|�۶��h������g�{�D�C���p[����o�B5e*����N��r�9$�P������N�]o�ޚq���E�.V�!�kU���:)��%�KgG�����/�m*��jN��:s����e��ރ|�r$�Y�@�����9�S�hN��CӖ��p>v��1�ɻd���5����ܖ&�˵%~���>��������/��LHk^�(E��_Y=J���񕟺Q��H�� %�?��U����J%y ګOgyo@9$�$}���؂��7vxA�����l��~^�`9M5�bw���>�=X�-�?�@�$��ʪ��+%QpT�9�_,�Y)X�+�j�̳DJ0-�ZÑiA;MeRsŭ\F�("%����࣍F@������b&��(�3x�P��U�ދ��h��&���Qks ����j��=�*7��?���o����k#��°i;n�*�$L�(D��st��{8Ŵ�"�<���4���n�sJ�=n�#�7�8�<��N�9�T)Pa��!�0��/D�d8��A?)�V��f&˽�[s�>V �]��>(+kz�y� �:=^7̳��a��B�U�;*����<�d����]���6a�:/���<�Z��������N.����[~r5�ό���y�>0=��ZC#_� �E0�v���#A�5��BU?�|��e�>�[zb�a�}��i}�+�'����:����t9)�����B
O���Ƭ]</��I_��8�d�0��y��èP'Aul�$
4��1}�d�Z��bQ��)��Ț��O��W�K�Ƣ����V�\쀓�B�CU�I���E�$��\�/�$කQ����E��,���e �`�����+{���AP�f%�/&���㴈S�8 ���&f-{�'c˫Dx�L2y	-D�HI��������O�������(6��. 5�Ϲ%�����uH���2���U���p�>ш�T��yw�h5����ˬ���5j\K��5����`B0��=���M�������U�(��l��/< ��g ��4�e������I�e�cَ4e�Ե��
�QoF�>T���u����_L�:�$���`�.ZP����m@��;�8j���<i=5�J�������'V��G�!���0��;�(�4i��;���D��Zn6����%W
��RLm�4�@r�@'���m�g�J��&�����tq�淹wѬ�Ǭ��n�� r����đzZT�Fr��[M�V\[u׾��to���8}4�H1��F�T8�@��2���: ?z���5�����<�_6��p>�F&Z��z�?ɽH�@��1P����{�����'�{�ĺ�F��d漴��L�G�D3_�a	5����ƦK�� ��d�{�}�A��mA�3�d��	��{o�vh�۱�0j+�e��@��ɠ�A����e��HG�}�� ����m�}���o���I�^��AY�ݻ�ɠ_�T	��,�;-�p�]j<:1��3Z�qc�W��i���z�sO{K;���|�+`v�N,�lu5X�!�ݿ��v'��.Y_�@��fy
h������	Ԁ?�u���==�������TRH�Y��N�����cۓ�$��<#A��+=�.��zoD�9�Q�����X3�mk-�P&��(i�B�-M�-���L��%���{l����Z>Wy3�ˮR|!���dQ��e��t�X��qs��Ǉ����Յ�h���Y�+��IɲB܁�9��W��.Q�X1���&5f^�2H�+�k#7��ꇎ�~ ��m1B���,�	1%�}�%��%�K��,$�*?�:�� ��+>����y��ƹ8?���]�]�F�L�Y��'�P4P�gM�C(�6�}c�:��P�� ��vd�
f+9Z��V3��]M �ܹ9�|�����-�\��fe��t<��$��5�:�y�
�Z(�gZbQ��E���X�ET���~'�[�&8|Ȗ������j�9Y��;GJ+(�3T��`9�cqjң&e�RI-3��56�H��$���Z���6���5n��a
�L��zp+�;OH~Tf�M�?�3O�\�A���^�BC#K������Gf�x��.0�~|-K�6R���1�������e�� ���_^��.���'�ҀG'�U���F6����Z��c5�b��i8}G�: =�"��O��ֽ�0s�)���˗4���u�UL���a��B�|���]J����|zh̑k���F�/�)B��	������y�M�E�F� �~7\�$��_i�+a֥]w5Նj�89�7��`�̲��tAn��+ �D8��N��:	�X��W�D]����|wj�KQ/-�,��KRܶ��#��1�_��,ݙ�;���K���P=�RL�KM̄�>�ʇ$}�t٠�l�Zm��0#1JA�"���������M�ld	��S��Q6m���lg�P�?��8�9��w3T['	z-�80>P��l�����Fmq��E��.S]�z�*�;G �=�1�u\Ǵ4GQ����� j�Ggr���h�anۮT���M��|B7c
/0�L��S|��r� kc�n�Mu�0�BU����X�sei�{�����Լ'�1��F�V�Ҽy��ʖf���� ��i=P��Ħ��HN���e�_�MG�@��ͦ��v��)�����AT�-�!���4����^�ы�T���i������Sz5��[��L��B��p�A8z��j
��*��P�Y��-�xX�T3�byݻà��5� ��;.����P����Q��5���SJM�]7�ͭ���s�+IĬ���eym3*L�9�>��ы���0�7���U�����C��<dr.��A{��
�NDs��\����D%���O�{��1?��<笧���M�v��^���^M<;�>h�.^_cGӴ��r��C�������~%v7��1�'a����'l�r�	�jf��p,E=k�D4�P�7�r8�ē&���VϞ[�G?I:����Ze�q�z�	_�3Xy�Ns<q�>j��b�( �Y��6w��࢈����H4��Fty0IƬʆ�����i4A��7!�#X�eƴG��z-H �b�f���햆�����D�ޓ�~�mc��Y��˖9,44�����.�*\EИ4���}��A�q�j�������)�}����JL$p��/A��o0ާ߮�Q"�\�7A׮z!G�	7��J��A�l�AE@���n�up��,��^��!I����܊�F�ws��r�[k/������ ��zJA�)NI�N��o6д����(��_��lo������6l�+�6�/fE�=-�ж�	�u�<�!-�.��x��s�ZHi6D���o��mQ�}8]p�#A����@��I�P0��2�3K3#��u$��ɪ�����V5~�/��t�W����q�!nzD�
ϭ&�@����I���J)6C�]5��]����գ��cWNP����],͟zl[W�/�,6�
5 	�@i�k~�m�S��^�j��K����jV��*M�$�0�4�R�:)���ٴ��Z��m��𤽳��f�~8�b1�Aw>5�u�4�(��gKbj��`'�C*�H��6!׵]Ǟ~�LQ����?�*͟ѡ�Z�t}a �De?͗a�9��E�+�-[&�<��sw�[m�^�s����S�u�� t8TpXP�+���'vH�7��������1+���U��0\U54J))�<+�s���z�(�M����r8���������fo(T���/�����I����ŀW(�O�������_&;L@P0���:kqޒ�
�e��d�rd�*hV�>���:1�'���n�>�c<8�U1�d��ޞ�؇4k�w�	!ț��U'��b;�ߥ��/�������|U��n\Ψ�G���o� n�B��ւ􈓣������lIMZ!�����'N2O���CK�4 �9A<~�
KC����|�mu�	�dHU����$$ﻱ���?{ݠΎ���1[G�}p�A@�D��-kV��f>�}�h�{߄�"��O���BJ��{�X��}��Aޗ��A����b2��Rƒl�Δ�� b�A�%>I�Z|��·��	��;a���j�� n���p������ ��:{E��Ν>}���i(��R	�$A�A.]Yh
ex�ɼa~�{>�jUWR��酩�X2�l��<g��г�%}ɾ.Q/��J���X���J<E�U���P�tU��e��`�4��-A��cQ@�@�&a�WpL9S9<��:N�*�k�-e����;�5�u9��-_�`��ge��'<nOw���

�x>`;�9t�R�N�/��[1d��S��*��oS2g7����玌ߝB#�U*��"�td��sSR�xGݎ���\�;�Oǭy��`���S����g"DaE�vl|TAA_�UV��x��#�J� �Kn����,��L-B���*R|�Im�T߲�z�dX��CMI��PxgD�0JY ~�:�{���}��AA�`�&Ǌ8�����sk�P���=H����	5���x�"��m���IG�yK�Nv���t��r�8�9dN�U�У�۠�����eK0!�7��X��!�O��+�5$�b�	Ͼ������P]5L�Z� o�QI�pR�w�]Hʦ�@*��<�(q Tв�06y?�����
����K7[��O�H�1}g�����YC^g���c�Q��֗>b��q�mQD	(hy�RwP	GXӋ�ӗ��� 2�Ш`�v�qU>+^m�67�d�>%m�e �݄�7�qf͒c �$���>c���]zE��v6�u��f�����š^��ɩ���x���^����~1�-�PW����H�Yp;��Oӽ��}I�k��9�1%�~��V�s�f߽Ǩ��@J��7X�:|m�ؽ�jH[coN���	�l��ȇMgV���<� ˃y�tq�1�hI[�{S�z��^j�?Ymȣ\��&;c&�k�q3����ww���B����Y%��[5��cE�Ć���BZ�P4�2w�AoB�J�G�O=Y�m@1p�%(�qAȤz\�=[l(��3���=7b��%�����ج�3���i.�'q� q�eۺ�@�e-~��X��c�\:��&f�\��Kr`n�O"�Pe��W7��wRd]�K�Kq9xm� �����
��3��D��~_D#X�I���`�"�i�����IU֝�J��������2�	�Q����w�M�Ykʙ����[L�:L0h9C�iq|7��?2�ٰ� t��㉭��@��f>$���k}cmx\ǉ���Ё�'t{����]���w�{/FKg����������{�ł��oxޏ��5d�̵��+i��4�֑�@َj D�y�4M՘2;�)�L}��;�q�8:&LTBN`��0����(�0?D
��-D�`��x�ֈs���D��R��[p���\�njt�\�^8��5�͌�)�=BN8��3=r=�(��F�U�)Od��M����Cm�`S>�r�Ծ���^_��
�,u��;���R�����+A���˒v�4X��ؕ�j���뜅���C��~�Da�Ng��Ԥ��\�ĭ���|�SE ��7
	��ѩl�Ho���lK�DS��^W�F�D���f"	}�Tk{��Ԭ��_!�U��ɵ��AD�*����He�:>����oNG�r��k�F�s�,�YU�Ī�H��ڧ�`��Wݧ�������˾�^��^���H��m^�R�iK��ߧ�|4zٓ[f%ΰ�'\:�NZH�B|�����:v�����V�ƫ
����uj�/�+c���A��-t�^q�~�A��RH�xv�#�|���1��"�����r���6p@�%<xz�`��~�(J���tb�L�>�ž@�6�3N�uf\d �Cr]2|�β�%T=�}��f�#9h���O[Q� �ɕ!��PD\
`��f��C~��r5���c$��n��2�FL�� ��7�oP̬9I�sޛ������.R�s��
b���y'^����l�����(]�+�H����(+M'��Z�������]�NU3u��dz�,�r��d���C�e���+/5TJ9�1d�9 4GV�����F��u�o�S�sD�Q�|kn�_��*��cW䐉�*�9B�($�1��̓FF"�=�\P��ZL1�z��t���a�|�zz��x?��
Cu��7���x2��=�#�U��--�|�sI J�ɔx�^OC~�(O*%�p�_N�-Vsw-Q���B�Ql�Js�#��U,�-G��[98�L��m�&4Y,kċD�I*�KNl��|�N�\M�J��̬�=�����M�6
��F�WR ��� ��#�43#[%����F~;�e�F��\����ҰS�#yu�)g:�wQrv��Rӟ�����P��`��"����$�ѝͣ��i��VVl7�$t</t�"��y�s��O��ɔ`)h��9��oHLp�pLG�%9)��9��Nu��W��/�%�~�|`<�?+���'`�~���s�{B�Ȼq��G�/��F�K�ѣ)�NS��i�;J���WV��-�&!�����,I��`#��(�*{	Bxn�=Ԝ�F��<��i!�K)�LY���&���n)S� t6��m��2B;��ƨXc_��}�.�j��E�[}�������5c�����  J��\���"/%����4���`��"��$��'�	�\�!�s�X֍Wr��U(A0TЍu���6Ւ��q��GA;d�8�(��d��r[>~�^���Ρ�ߣ�zij2���o����77/M������NTH�)i��T��܂�`��	BIH�DE�2�o1�;�8��;+���e�YsV�k��VAߣ��.���P�7��5���kmxÙ��&]�j%��u�d(��z��&�������H��*�k����N{\��F��)�o�V���S4
Rܾgb j�d�=e�
i�䬳�HN5������M5gRe)�"-��D������n`Se�C��t��v�S�?�J��~UmCϾ�M��l�=j�oz
�:P��U��~x���W^��:��1��x&��W�S;���N,|d��3@O���h���E�"/�@.�S�j x����ʃ6��Tl�{=�Ȣf0]���8[Ep�y�8�X~8%w�!QRڱ�n�a�[$��0'JtG
����Q�]�F
�$��@�)*|o��͓������1�b� �}��g0��qTf�8�)g�������R)3�1%��Z�;S[Aܔ{���r���٢�'����dRd�
��0�2v��f�#.:=st�<�����C�2?�MW�m`�����^�G��Eڀ���$qق.���Ɏ�?r�ӓ?;�Hd	t�	~(�����X�plZ|̼�Y�=������k��"�#�ݮ�g��Hlkls$���$�]5���X�q-�cw"��7+�܁����Lr(`�B�qW:�D1jv)�6�Ny6��j�g=`�a��L�C@� ��ܦƳ�(,��[����+`�{H�����IR���PA���Wc2���O9��E��(�y� �O��˅�C"K��5��.A�V���\�čc�l]�A�7�s�g�N8p����\���k�d��~�9���i�������4��&��dֻ�d���q�l�Έ2�ĜNfqJ�JU��R1K1���K�[x�y�-�>��k7p��.�_�aݔCO�i����P���+���L~���á�Jt�7�?ϣ���f����>F�x8�=^�:b��,�St�q���Q�Q��I���Kҷ�
���h���>��ڪǓ����jB^N�Ԕ�k�,�����)�/f�[8wa��k) %w�m�F����X�m�B���0���|�g-��!̶c��%��(WO�?�ji���{�f����C��<�fJ
��\m�#��dS�PK��JGHA����Is�Rn�Ch��6��*�CCs��|%/b�)�[�gDm�J�q������[2s0������q�H�~�A��ߩh������4��+����M�l�5sOGr�p#;���=�BO�c����b��X��B���/�-,.e�ٟ���	(=�
��~3�q	�L:!��/�_Q�bHB�W�%[\�S�>�<���2�" ��we��l%w����v`<�> �C>��%�b|7{�tz�V���7��T���������������`�j�Κ�	#�mѻ�����ۖ"m}4$J���"�M�й�u���4p���>Y�xW����l��n��e�KK;^c1H���'�U���y��2p�<���A|0���O1t��tO6p'Sb�;�f��۳�MМ���0��|P>!s��6w-k��:݆�,n+����H��UO�׆"�};����;g��=�V�i�ʵ��]0K}&M�H!��&�#�$Q�$���|�$ >qL��4b�W�b�#
���WG�!��a��n���X��>��k)5x:@+�w,gH�A�6qaE��jl,E�z��ĳ���;�����l�JP�qHꆲY�e��˻H��"�0хGo J�hX�Wy+�b�h >�6����V�;sB�]Y c�L�bO��)�t<6hl�k�ؠ�(�E/�h�&LB"�������N��x�>�U���������|�Z�X�(�mvj�n� ��]b\K:*�j?�!=2��ۯ�[�Pp��=����r�O�c�/c��,jltFB���i1���y*j�n��j���\��(�TnpO����7��N�o�<�Ըe�����R b�t�<g�r�C�s���R%�sζ�n^��,D�j!�~�ϛ�AG���~(wr����⯧�Lǟ ���@QU�4��'���@b�}��i��̫o��_D�O*w]��N��>=L��NFc��h��fz�[c���uZ��"��1}����Nn��(J���ĕ��A���	�2�����;t�(��@���r�ΊLA��c�/R�Ltlwk�h�C�8�?��=�]��>[o�j.�X��Nl�	p,@�q���>:�v���w<�w~��PŢ��zxAdVr����;�EX��S�8�5^��o��\x��▣#���aa���Ikv�0ΙP���/k�KYʭ��2k��Y�J^	��L SS$�7
"�?�D�Y��M�+JXM���	��6���������e9gȃ��r��&������r��k�f��z����,|��7rBٟ�y�w�oĪy�||���벽�S��{P�1���*p�u3[����ۣ�#3�|��-���@���r1�(eC��v��<�< ^��U�xւ�Khܭ�_�:���.���,���{Tjp��+���\�rajd�K��C��pd��*	*#�{��Y٪I������I/��NҮ�-��XFѦ��d���]T���ݑ�g����R''��) ���6�An��j�w����m���E�2��1ptNdS�f�˺B �x%��5�R�!˜-?����CU�����1����~N�/�N�Xe���'��},<���v��˻q��`���{��	M�mH��q���ˆ�ދ<�>�!���k��^]-p[qT�%#�'q�v���C�����G$0���V
�	O�ku/�����~���2�"(�R؇i�W�-y@m�҆l)X���hX'�|F9&����$��%Hy;���J���|�V��V_��4��m-I�n�T,p����B�GL�ó�A��Vi*��fMZ��T J��O[�͈
3e;Y�����ۭ��r]eȻ�4^e�N��	�+��� �h�Z�L)?�tY6�&&�j��u,+�R[��pu�P����5\���>�
=[u7�.�Ѻ3�~�4o�u/�W�"���!����`��"���1��X�oa�z�'��`1ꪡ�5<�$�MP�)�׍�h1�+r��������)*�\�=8;�֯��>k�r���Ky2g�oǝhkZs&�e�k'H�T�f�Y��ߍΡ,����WB���g��=y�%�l�i��yq\�/'X My��Y:H��u@"�Z!���j;�� �th�� �L/�0����/��Ec��e~���P��xo���Y~�]���:�7�>�CO*B�&��x4��3�жnʾ�_��y��i�����d�����X/���$Y�LD��u�Rl -ŏ��Ӟ��<)9(B�/���㩎e	�^��F]+���\���|��_���ӌZ��X�M�����C��?z_�� l��a��x���)�-�X�j�n�R� Ү�5�GE,�4~��̓s�g���MW��0i#7��&p膡������m�y1q#�I��kj��c��I�ƺi�`�u��,�ł!i���#��ϼCb#d�w"�����b�Yd���ذP$`�Y��6�HH���J_�q��|���S����Ŵ�$��]���&��u����Y���3�s�؁%����&К��Q��i�j�/�������&���`�:��OH�u��W�b3;��T��.��A���u�y���9. �����p�	����x�IF�pH��@	�5��G�VM����V"`���^^�q��1�ۀ��>LӣC�Pb�R�����<Ѻ�?k������K�~�(�c����G���4n L	|�X/�:҄�WJ��=���3F�X��G��kϷc�/��Azk9��>�� vlr��5�B�h7 ���^�E�����gz6�6V����t�婆}�ی�t/˨�#JS��_X����|_�� �0�C�F�Vm��Mr�5?Wʶ��.���H��4\���i&v+y�X+N�}�i�x#D��'�"��/���6
��۫t���	_�Hb�O3��^�g���۹;Xg��۸�4�<���Z�xXjL`�}�UH�Yf��zr���w�\�\�/X�k����ɱ���t���V^v���z�x��F���DȎ�>�'d�Z��\�Y^L���s.�riv�n����#+p{m�Kg@�D�U%���El�"l�I�<�f���o=��af��sB���cJ���՗~�o�ߎO3;�	�@�H-�U�_d��� �#�-���`ܥb2�gK��xt����4RF�}u��㌫5�u��O{�u�@���d��2�.Q/�ֱ����@&��*���U_�_�7m������p�?�=�����i��A�T�+왎u>���R�LGC��˸y��*����㕑n��^�]O�W�
�s��g�=t�B�_�v<d7�3�%�iY]6�8h�oџ}�����l'����������hm�A�<�^�}�R��oD@�r�����=����Ko�"W֜�Lùw�r�w]�U�]�_d���&�4�}['F�Vv�/�táG;^a�@��}��<w��V����y�t���Q���$�`N(�6�M<�"���3^c��[):��/�!+�fFx=�u�>�yݭnL�'^���)�����_���t�N��{p``M�G�I=��������� }�{������h�R�o~y��"b�>���A���p�V@|��F�ӳ�3T^V��쳟�s�]ڄR�-Kv��󰪤�����nCݒ>k�k9"�r�=@~�X���Wd��y�T�ի0��1�+!��v���l��/h/�Rn�>f�
���b��}<�v�i����ܞ�W,�����<��W�1dӬO�h`�pq����\�tk������s)���+�f}��pu�-�Cx��WPy ��J�� ���RQ5�lfȣ����S�S�+|��&8���������[�k�z�Ǳ������NKa�O=�Gd���K][L���t �H�g��Kӑ��H���&iF<��KT��4���/Au|O�-B��?�`]�.Q��$���ύ��ҋ����;���2��C{����}Ynw�I�_ -z��3Z�(�&��j�Z���D����*j��W���/��I�׼,%݌d���)c-���TlANǺ�Х�PV�o��N�bT�ߑ�P����w�vﺟ�n�],����I��6�s؀{�\��*nU���B��:�'~�k\���l��*�~����f6���뺞F��'�{$��E���2��t����_�iBumث��]��IqWlȸ
k!;���D��c�q\vu���aNW��\��-jŎC�"|�n�M.TY�����y�T�=Ɔ�h�ke�N#~�\�1��l��醝%4������IQoD��+�ѭ�,\�Ǚ��yϜ��_�@�ԓ,A��Œ0q�1`�s���.S������-0�O2`�<��)��䵪�p@�eP*;Y���'/^�4��m?��z�K� qu��P�4>��a�(�!Pu�c=o!`�ʖ��p*�
�����H���z+e��l�m���U�8 ��I�c�֟��9�����V�p���#A��|̰m���>$�aᑳ�U,�Vp\0���P��|�v�޾�٘	��0"�?���ˤ�KoO��;Q�Ӓ�?y��F0��;Վ`�Βv�k�7�{��!��mS �:�Ͱ^�Y�z��m�|�3Q��͞��Z�D�V?k�vQ����%MJ ��Y���؂C'�x$'�W�r4�莇��'ˤ0[z�z1>y���j��:zH��٭D�}{h\��5�a���tES�,f�%�\��z"U�@Lt�>���a����iu�����<�r�����-��e]� q�µO�O;�Ф��v���&/aB��w�^w����.�-��3/�oR��N����l��/BPZփ [ꐼ� �;�*׆^ݰ����_ ����׶��m1��L��08
��"�l�+Ӻې~]��%�E�y�|�#'�yI��%8i@+�㞧U#�n��.��w)�u]@q�Q��2A���~�e^��k/~8��#�f}zzv��nc�9�Xv<7s@�W��$m�o����҂��s�.�D���f��n�<�F�r�p�ɝ�� x*�Q�8���Q���-�j�X�5dح����=�p텄XVJI�6�Fq�NW��((�MD�����J��n~��@�λO W�"����-ڼj~�@碙HQ�|b��@�擫�R0Pݓ�07_3N_HYf��7��Mc�x=ji�mR��/��u�tќlP���ͳ������9��a0c�N�U���gE)Pf+>&:](5|C0��<�w����Q����u����(�����T����F�Y�dM$�9��Ԭ42F����T���6����1z��6�PJ��4�_� �s	/g�]J�-���,��BZ���$;��R�bp@�ɫ��i�k��td?�5ȥ�^Y�!ǚr��Z3���H/�C0u�@/����{��c6Xu(>X�%ݾ&d9�9��1����rx��J5%_ӱ��CN�B���AVb5�d�ǔϳW,�HS�pL(�\�CʓaZ��� ��d0{}���{�Zg<���7�"�ŷ��d�f"�������]7
S�c�\4�RC�@I���Ȑ�U��G@1u�$4�������h9���s�}� ���=���u}t�"iqT�J�c[2���K�l����vCm� m�W�_�K(�?��D�`E\�QC�u��KЉ�A�?�3���,\-י �v�t��qؑ��% t���o/��L����yM�`��S��VaG~Dg��C�F��t0ڥvBd�=W �Q�Q�ȱWퟞ�q��^���(�V7������]�/�錄98l]����9h�g�P��i|���0�k������H��1e�=ޔ����,���o����p~��F��)H��rt2�f��������S�5�Ӈgn8Ũ�C~��kZȕ�����r�vmh�o�-��x}�9F~�g�C�� ܍��r>����^
R��Q����h�u�d ����xN�xu����'��ϙ�]Ky��_����+����J-d�~��b�db�r�b��Q�}Lј�-���!�b $�Y�~�h5�z^�!�����@��!��I>#qq�g1>D�52^@�q��k�7	ϦX��+R�~2=�H��(�8���@z��W���qQ��Gj�C�������/[`����s�S.�����I|�F�`M��1�ދ�+����҂(ɊH�J�V�tW,ʆ	2�^{�h�"�����G�΢*��)}*byqL �x��C
�e��y�8[ł��k�M!NCQ�� ْ�q/����3F�����]B�eÕ§r���:`X�o��K�/D�u�X��S�p������*�i6�6YjT��h���?�\�Xd��(�,?^��*�GlCs��c�C΢�qXy��Ħ*K?[.�`��.������L<�eU$���U�������tʌ�݊�'���ϐ�������Y�T�r�βң&�7u4�(�5�]� �����M.|7���ǣ�[� �ԦE�M��k�I^ir%�c?�iڎ��B%�Ĕ�^����x���rE_�7�,�|�7H�&�]���P��"���W��,,,�g������,3P����.��|0�eѰu0杯��y��5(�����jbW�$i� G^�U*���"@~	�ĺf �+Ə�e����I�R�X��|%�c��h]z��~�f�l��^�W>�����NN��Ee��p�ѥq}R�񰙰�\d��X��M� Aw�d����(�~��L9�C�#��,B��ε*8��k��AǱ��`dr��e_�d��2L�ϫ�j��tIm_*F�I���c*�U���a.��Ѿg�*A���9_U��8"�lK;]��ܻ�6����bb&��shř��,1i &w$����{7�e.������1c����<���� �D˧�/��ջ1�y,�U�Na��T�`����R���<�VTD>#��.<����LWr�]��"�	"��)">a����l.b�^I�\�	3�K�klGmBI�f��f���9�Iѻ��芒�Ε�ː�q��`��[ͱ�E:)ZU�P5W�٦P�ɫ���ԃ5�ΘL�]������i���P��O�k:�tlP��Һ�g-T�mh��F��f_�5�J [m̓�X���eB8�j�ڨ�����Q|���/G3޸̛g�f�J5�����SR=��}N1��d���殭���/�ovǚ�	ja&x^�;�
Z���@u"�O0侊������Nݟ-���@7U���%��8��� �#Zxa��t�8b[
��;w RS�N�i�X~$=��l�x�x�������� ������C��8o��0�V��+g,�^�����C�	�k֪�k&I���\<��i�4�4!��<E���`��d\t�{c������� Y��^Ҍ�p���)�.ҴN��ǔ*
�x�:��h؉ ���w	���N���J�r�hi����H�<�s�\r:�i����%٠p�p�Ѩ���?�o\���%��*>��q��3"���i�v��!��m�N�)E�4���V,x��G���u�7 0�`��#�D]`�GH��\jΌ��.�2�l@6��3�'<|w��Cy��׍����*�D�E������09E$��s���-Iq�����B�xe/Y�`p���^���M8�qS��j�ZO�[�h����
P�;wQ(F䝁9�#��E${>�ن^�X�EWS�2G���kTM�����hJ�.(��c�ZHos'p�##��	�]MYm^���o#~���.4���£����hlP��[|t5�h:�	@�]F���s�o���v�F8�Iy�p#��8�e���\5o��X��A��M�s��V�2�6x���(���,,w�]�����������}9����@5��/�d�J	�����a��8]R|���q�e��3�Fa1�T�cS�_L#�|����w���qb8�9���/:AyA����5�-�m�>�ۓ;�C�}~bׯ���H��$��j����X�b��\��G�����p���i�햫ߵɎ]No��1�E��}XŔ�#���19���p�d,�3vqh<i�JȽ���ˣ��d�������={ �uу��A�.ɴS��C�J�|a���G�Kn�XN�����Ա���[�=�,�Il�D�ڎ:P��i�T�.���M����N=hI��� ?[��Yη����)��ﳖ{�[���h$|�EB��S"1��-S
�������gI(��H��B��>�7����׭6�7�d�U�>yKi�B��^��v��W���^�¤���+�@w���u͝E�߆P���v$�SzJ\�!��5C�x�̸\.�W�$xP��:�̮�����W x�c	[Ihy0WGH�W�&����=�JE�I6 A����Mc��Op��[���|V% ���i��Z�o�g%��hc}�K�~���R�Z\�����/jT��b����oF��߇�q�ײ�/
�`�Wa�M3����������1��]"5���q?P���XܗF�D�d	H��č�����?��|�j�QNIR�pHq������"�ב�;4���w|�lN��X����E`���m��1�����ͯ�W���K�f\��S�`6)�&���+��NѮZ}����&�)%׸����{-8�.f�G��'�iG[��R�+gr@��g\[[��������P)�����e�Y���,Z������	P�a���^�o�
�Kp�z�[-h�Q���#(-:)����Ѝ+��WkQ�3Ri����тQ-��8�D����?�00���gVJ����4O�ms�&��i��N*��==�u�g�u4�DN�(E7��|-X�Z1$�і����\��k�;�Fe� q?�����/�����C�6n]�CdE$I��/5�jC��G�^�*3�	{�Y���X�#X�`J�g��3,e^ݮT�{ʖ $��O��~�"�#
��Mh��&F���L�P˞@	��)�j�8������cH�Z���J*7��Ѐ���8�$��)Cţ�l�����=��Ds�������N�bO�E.��I�Yל�X�b�
�����5���a|�=m{"�?���5�z�TM����ek��8�� ���k�@�RB����Z�N�A�w#,����;���f���p[iD�.Mf���F��\2����@�*gʘ�K/P"Oh�׳�3�İh8��O���*��	�Ī��f��~r䈽��U�%a�{��@��J7�>��<�+�p�#�f��=�P���[HaC�01��UO��x��J�'ړP���ՃZ�� ���4ɋ-��n��I�m���*�҅ �8y����d�y��N�FP�����}- Gf-Y�����!��S�p��d6}�U���H�LhE͑נ����E���&H��H�?�Y�ܰ������D�a���v3�D!�F#6�je��d��Դx���J��ɻ�p�7${�x�ӎ�]<�>	�G�ʈ{7FdV�P�H��*�{�_۫c��K�ze,yw��0�/jH�6���:�b�jf�ip#�/|Զ[��S�t4���˺���aW���ZERid���bvG=�3�7�2+$�g\/ձ�|D�iɃ`���Ҥ@N��U{��G�b
&�a�g?�~z)^�`�x�s�`���}C"q�A1���Gyg��r�M'8:X�-�u�nʞ��Y��{D�_��ֱ��ͣ�%1���7��#��#J�CN��"��l�V�T�v9��Ҧ�o�������
��N ]U�7�+)�狚��J{?��t�{�R0�Z����M�$�������[#>�Z�s_Y��6IH؉��Q��! V��,=���m�J<T����Th��M�
����4�����`����GߧӃ�����b1�1;�������H�:	(�=X�m���m����6@4
�.5�:Z�Y��'���vm�� xK��<��-;�8%�IT�폕���3.e���s�x����ե֣�m�f;:7��M���������c`��qx�g��k�`�v��By��J�w���:��&��0�� �U�P�Aa�2��6Ô�j�z' 6��@Wl��u�8��4�3���˲W�?�hl�djK.�/I�?�����J�5���!�+������~�K��܎M���7��$l�r�+P-��qn-��LQda�`���/������&
�`�NI��[W����<PW�ؿ��O�=��I�	}\�H��S���̝�}��핼�]����v�4w�I;��5�oM��t<Am'MD:"H�>U/�f��m�A�ShO�������N����>��Z�Z�����m�Y�9=&���Bi ���|]���E'L;��~d���js�m�)�ҟ U�.�>�xl��X��PZ��� ���L�pΥ�1������JR盄I$xa�#6"����@AY��a�9��I�/I�J�����'�]�:o��#�H3!�6Vg���o`��g���^�~�3Dd6��@ܻ��m�w�<O��]n	1Ҁ����֙�n�a0�����O�F^�tDW0�S��B�.�x�N�Њ�?w�J��o(��� :���"w@'�	��sȗ�?i��8�X��2����A�e��v���h8E�q�&�O×��N�r;�<�G��M¨뫨�$4��Lm:G����+��w�3���P�G�8�wb��%q�ِ`~�v�#�]���7�&�(,{_99r�U�g�U߱�T�����#qH�8`��:��aJb�qB��q�w�{J�P�j��UD
em�`��B_��/���.l~�\�T��	6E�N�:�X�3���`����tD��a��0ƅ��Z��/��FE]Is������f&a�1D���4]����6la�g(ۊ��B%-��oL\9�������}B�D��P�٥X�/-�j�2l 3�6��M�C�.�_��je���=�����0����Y9e��cz�զ�'`��*f�.�� ƶ�f�
Ǖ2���^������:s��q�6#. o
M?��F\�_| -c�}
*cW��c��h��^�K�k˓(���s��M;�[{�w�^���,����H�,���]��b,�e�%���ʥ��Yc�߬{���CS�Ɵ����>�9�</2{�B��g]C�k-�W�?q�H�e��|ߵF���v�f�$Dԡ�D���x����}a~�����0tJs���wb	{��D/}��lE@��������%(O��hD��vLEn|.��|I����$���A@{�X�<��h	�_���|mF^�6��:x�D�4�O嚹|�����4\�H]�8A�6�*z�TR���uL�`f��<�i�1�'�K��~�T7����%�(Β�-Me0+�Zb�-�UNz빈dE��`b�{V1a�y�4I��X+cω/,
�A	��&���V�g�`�>C��Ap��wz�a!Z>�|ڭ�x+�
H9^�f|��E�^:�xж���j<5�	]�	����
}x���0�mE@67
Z�n�<�߬� W5��1
a�e��,@�:�r~��w���.�V�6	�M�?��dbdi[��(�g�z��d=)k���hI��,+o�K���Zp�9ّ�aa&�I?�⣱���ϝ�!m1{���
s�~-�鐜�������ud�4�F���Ӵ���*���PܹW�����`���Y�[ �7���T�sh�/���A�>Н~�Y�ʋ�J+��}��F�9�_c�ӆ�U�e��
�n2ҫC��_�\���U`��ij�q����=�$*՜���0"�o��]镔R�ND��;���f�"�����3����V�d�u��DKq���:�иY���<�ӸG[	�
@�p�g�$M�Z��Z·�ιgL%�4�k���B9 U����9��gQ[��D.~u_/�]J�Æ��-��҇˸���LL^@�����\+}��d?`O���>^g�*t $�(/������&�s��|c��f�z��!���∹����^q�

�Vl�\��Pyei>�f�^�Hϰ���}�(w76�<�J�n�X;�h4�� M��{��ke!�3�مM�<���0żlm�p���'�Y2v�\�4���d<mXf^`�_Z�j��<����%�:P�5#����l�5p�E�M�o
����.�
b���P���V����H�i�� �Q��%���f�ȑ���s�W#w�cVm#��ܝ�Bw���1�*�7����c�۪�U3��R:[�Fd7~�]>&��^Aڧ�Q^�f�,nU�|G�h|�mL�l���A�A,Yk�r浭:��J9=�+��1#�f+�[IG;o��u:�fk4P�S��j v�q��	���N�z�6T�? ���Z}U�"�̯����7�y���g5ʗ{|^P�(��H ��ĉ?A4�Kjqk��r~��	,��-^ 6��,�)p�M��ފ}�Sa\V`��Fr|I?���@�>ݧ�D�8�u�E+G*�h}z���m�80�1dR�r����3�I�|p`��Ĉ��"Dc��<L�Yȡ���%4�!b5���ȗ�\"��OT�_�������F�?�[ѳ�����z'�(��7n���v$&�s��	��մ �G����nc�eb����#��G8@$�+Ʋ�!)W̗�ǋ*�dԘ��J��៵�~�h�Ns�� ���k��I,�S�D*i#N�E�`�a�y�{czPa�h������[�K�����l&��Yt���nBN��VCu煄�Jా�<ĉ[{���"d$`��K�/�d{T@fx��*]�e�r�,�*�O����J&�_�nR��mN��d%"���i�*���]�4����		S����`�}8�<����!��R͠�Xc7�� �+6Pt``����n�'����hf��#j6Z`�M�o����i�y�.}��S��$��c�YZ�_����F�N��Z�O�*�Q`
�����
�Ќ��(b~͗b��ִ0b��]�6ZewS��E:�߱{d	iI����GD�~!؀:�<?��9��7�ř�1 L��U(��!��H�?�c�3����� <�_ݹ���o�O�T�q:�{5f�/�+��F>���8�2���m������0N� I��x�<F�\t!0�'�'�֟t^0H�cO%��,ħV�|�~S�5
��E�Js�7C� ��|�X_GM�f-����{���BK���W'������3�N[��xL�{6���:�`�b#�I�����Qx�Kp�c)'�Ƃ����d������|�� a�D���oUײ��i�R��1�n���,� b�J08���7Ʈ�����j�X��9M��5D��-���2,�^���
wPr@Y�;)��E�fD4O^��V�W���J�qE�i��!�7�J�:�?ǱV�9׫� ���B�d�Nn�ec�Q�LD�A�k;�-:�^�y��/ͼ�
���'��o9�P��B��g)٬�G��;�%uk��.�f�;�w"N���.2�h=��n>r50�g�#
M7=�h�`g��ܤ�<�x���-��~4������h��$p�B?�?�5i�pnᔡf֧��>�G��<ļ�ƶ��G#�w�|���&�gu[��@��k$�!@�D��*�h������p��xp/�B���ז+;�"L����C�0@�˞
���F���z�1ɶ���P���S~�����ʘYg�����9��q��z7l(
] -�ڨ0t����tԲ�	�����i��V��y:t�ʢ�JQ�i��zQv�^���<G��'첑��~�i���7I�?r*�t��u����\��͛W!1c~�qe�S��&����?��x��aLN���TT71&��A�X�����	(��AK��$FQU/���h�
~�J���ER`���(�K��#ŧ,7S5�������6u?2\4�T�Gx.�DN�iR���(���i��5;=�*A#��}��nY�2"��I�<E\��,u��{_�٥W`l�j�����D9o�~����v��E�>*|Y��'O�l��椱������vR&-5:�0��W��7��yEQ��S&���C<�����)�����Λ��&�N'J�D
��*������W�����8ȩ��>+%���N��è�W��Zh@*���r�F����0i���G��z��0-�ݜ=-���x�� [�UC��SnhOz��[���
�ڊΗ0���k[ �%f�te,q��i'��x�Z��<e�yHNYfO*�"����a�	��_�H՞$�N��L�v��]=�Z���_���`#	M���e�e�G��I����>D�o���7��L���[�}ֈ��k[�>���k+I&�z�X��9:���f���i/�O(Vu����un )�RQ���\/�`�͹�A�E�Ç�ð���h£oq?���<�����LE��|��I�-��[��T�'��ٌx�Y:�9	lS��У?�є7���-�]��� ��5PAf\"`X}�~�W��%w�2�R���.�駸���97�R��b��.��rQY䛛�`{����-�?`�h������Q�ʦr�δ0A�5k��S��9ZK�˥�Ϥ֥u,Bӧ�!��s����t�Х�w�Bj����J���M�ͅ��f�^��уӏ/FЊZ�;��k/�
cW�ru[�����kچh�	"~<�9��-t��)8 �\�˺�L#��su@�~�ŝ8�Q��sͰ�Ѵ��:i�X�Qp(w�1�����V�7�k�ʧ��f�ۊe��0��U�������[�o���g/|��`2�LPG̞�3�A@ß���N#���4��n)Փ���Z�Q,�At��6h9~r�^��J��q�p&�p{75����c�yc��Pa.�����%%��J�,�n7#B��q��z�+��]�����˸I�صS�M֭᭧�w�bl�^����ܢQ��eC�5״M��*:/s>��:���)��V �\�(�=����Fk+D� ��{����Og�:�P�,~�I`RQ/+��h�y� )Ȇ��B`�Љ�}����n�����z$�&��j�_�5z�j֭KU�[������lD�ƻ�Ș�z�s����%��w��'�68i���b��n�X<�X��(vj�]*1pȆvBh-��Y`3�oӦ�`nʄ��T3��a'P~=�֚��"=�"�$��O�Vg<�4p��b��⨴D)��"����Ψ*q��"�0�� ��	���>�ώ���=��(�g�#�� ��P���KJV��C��#��pY��P������cՈ9Ev[����B������"���o��p�(��"������e�wM��cq�O��Td�#'�Wӱ�7�4o-��S;��&`�c�������~s @z�"������0L��1�*�"�T��	��5�z��Ʀ#��WΔ1"A8Pe�����RX�q!�*\���[����).F?j����U�|���0g����N�,M��cF _���Mt��̠���k�����ORu�g� ��`��t�:W�[���H�k�7�.R��F�m�+~+���k���9���:�`�<-ں8}��d��1���6�-/z�����;P����n�a'��ّ��O�u��6�r��{,c�^=>ܼR�z1�By9I�����IǄu�hT:���{�V��q#`�B�[{���	o\���G��ÁipR��__2��<�T&���N_6eܴ�uS���y��}ii5ui���t�>J��;a�\ޟ@�hi�z̄�� �\���6�N�o�|\���k���k�ף��G
_�,��[G���ɲ���%��kU{���h
�Xg���]���"��Op�c��in'�U���+�$倶� �,7无g�3�K�S��8A�
\��g����y-قg*؄�l�&a�u��Mi����Gν��6S
LV�|0f%Yk�ٻ�kV�#����8h��_Z�r�U��:A�(2�kd$����c�����eX)�쇍�����2��d?C����3( �S1�{�ԭ���~�W���o���d�B{ƥr��%��z�Sk!L>EU�~����P�:�߇��=���5��*��,va"��}h.U_�(��S`�M�.i��ǌ۬ț�,�`0��i/��(��ڠ�ݼ������D.��п���"c2�
�L�!<Q����iKZ�1f����)���c��Nu)��E��0�*�R����xk���j��D}���	ky=�#���j��Қ~���I�﫝H��j���LB�
WG�Dɕ�|^�p�q��%�|��'��-nEC�х�o��'��`7r��ljlª,n���L���Q���,�@���0tj����Ȃ�up�}���~�hq����'�L3�U��j�̟7�گ/@�}����8G)X)}n���wR��=$���DФJ������-\�o�s��.�vJ;�Fڊܞ�����=�y��oS��П��E�!�ٸZ$�U9�ͼl"�����%����j���"X� ��qU������a��\�ŭ�� �qr)L=��m:ff��T,a��m�QPOמ�䂗���Y;�� Ǻ9���K�����l|>��� ���1������������e�SI�~i�����ȕ[*��Ϊ3>�*2m�L�m��iz�=2i��i�[����h� /
~(���]�c��4�&Ay�zvش�~Ǭ޷�����M�04/g��X�� x �_I��۳���ķuA*fv��;H~��DIX ��e�_UOTl=]!�����s&k����&x��p��80���w����ϓ����U�W����a;jg]�k�e����_�����`�ZG�v�bF-/��8ט�\>xܲ�E^J�NsP@��X ���!�Xu���a��`�0i��Ƶt`��sέ&X�W����@io�J�^f%����䳺����$ğg��p/E�6�Fm�D������|,�EӶ�k���P/�>�s�ҩ�$��"�l4���B%'�I@x�(R$��E�;y?�LJ$~3�Y	����&�B�t9]w�U���\���K�Ʃ���&� EG��^;;�lUi�4�<���� �gmë��gJ�<�d������8ݨkffb��QL��,���(�"��a ���]wI7��v��!�>U/n0h����1S~�Q�UC�M�¢���T}��J����t a�!�Jq^U60�	kĒ��O��m��va&�	�<�c��'5oV�Q﯅��И�FTF%��iIQh1C�
���?2�M
5����)�]�5���*�/��?�V������E*��FQY��~�a�>�|�������yEzs���+6�?Q\"�k��a8����EYo$�4���г�&ߎ����0p��۠�^����J�2~�%�qq��7��K�~FkN	�5o�|�F��[�&���ӡ��uss�=%%�+�Kq�2T=�i�K���om�dUպ�s��~(q�}�p���Y"���+G��	d- �;�S�����[JUe�u�ʒ��y�M����)�8_;y��5;�B^�n�΢MI
[e�zɷ0v��et��)�fq��)�D�aI��S��������,��(�I	p혪��J���l��O����<f)D��2���;���-������Qɇ���k���|$`צ���s~xӁ?�D�6&����^@*Rٹ; &�g(�՘�x��՚ED�5��Z�0MN�|�z儧�.���+w���]��%�c�(�����$[J�3��J(�<	ܗ�*Ӛ�~:L|g��]�@e{yS,v�(�%&�T풡��x/���XGw������xT�e��|�ŗP�>�Y�a����7<���~�E8!x�S����SK7sb�qSZ����!&t��惫|7H��,��t�0�3���6��w��c�S����C�s�C��2� ��i 'M�o��3IЯ��&��/8\�G�E�I�3�h���䀛�OO�*<Vcj�`��,�-|�Wo�<�w�{�&uI��2�&]z.�-)� o�P#KH��n����JW�R==����Ӹ�	K��˨��H�2#���ߓ.�@Sďq9ñ%Jvs��z�;R<��q���ϕ�'�(�g��E���VϣYX���I��PIxZaiHU|3"t�ܦ�L�gSlZ�p�����a6�����~ d'
�
'X:�0*�=�a�Ĺ\�C'����#Zߥ�V�;_J���Ȯ8#�VԣŶ���[��v�����w� L�j����;|\�{��5�n�dF�s�OUT,�}�TK-ꔌi��C��}֦t��Ԑ�g:8�^P�T�~�̣����c���>Mzj�w.�9���z�d��EZZ�iH��ʙ���I*�� �6e�񜕵a�(�&Ke8oԴ{[�RQDj�����C�owq#zEA�[�RY���a���
�q�=8�8�Nf���|l1���8�*��q�h�#+��i���Km��	���oZ&��^���K�K�84������澣	J��#贤��Cr�$qwf�ˏ�`0�#�}�����w�
@\]T8����p�X�>§%�Ղ=�N��h�t*u�4����k�6e�Ȥ�����a?}�>	JOE�w��y"I�]�r��;"�HS
�}�Q^ƚ�{p���\�����u�U��%��^`�X�Z���F��ةE	9�z��Rэyx���}BF�v�RvB���]��Eڭ.].x�T�s:�0��2=%\fh&I�>�D��aG���juw�QT��T77d2!�q��_��<{�Ǽ*���G(haS)D3�ۦ(?e�i	�8CQ:/�"Q����n�A�~o��I<F�RS,�p���+��f�vL]PZ<�]Ժ����E���
���ǯ��)�q�#^ԩ�l���S=���<���g��ާ� �0;%jYt!�
v;���� �&O`�b�;��l�h]9,p�����><��f,V0��������1��Mo���n�e���c�3���L-ꆬ{��4T��g���d)��-L���<AMcq�0���\An�4�o�遯�U;������/_5�Ѻ��Z��b�ͱ_��LZ~���W�#��q�)�������qR����js�~�S޸7^��Q���%����E��!a(nq}��"鼧Or��x�	��v�m>3w�P~ �ѱ�'�)�f[5�a���	�Z\��YR�5�������<�s��I��oI�=R)�u�Ш���d����k�,��"ʛ5v����z��X�2��_l����|kg�	F�Di��P�ݕ`e�>C_ʎ^����(�� �~oo�*8��Y�:�+G�Y�r}�ݘd��9:��i�5�|,��f?���轺���Zm�k�w?y�{ym�C�I~��Kt��7&���~w�5/ӟ�Hֿ�x� ��ݛ`b��I{jB�7���'T�LsG�px��7�jbv�W�@6N<<���5ZA��?+��딃d�J�1�y��p��΀��Y��uc-��,��9�:Qt9�n�= ��M�kyѝ�?��%L�"��a6��M����7%X��Q�[�b�7q��)��ශ��>��Ɗ�ǲ�?�w���o ��C*2��8���X[�?���W�:W 6����n�� wF+Ib�%�5W�Ni��Q|�k�E;_�xk�A�j�~1��SB3��~�K-J3�����|ط���ѷ�>���;/��1#��̚A��7�����I�?@&x����>�lx��y��� ^Œ7�^���)6��}wF�}������-uf�������q��ZzP��C$��0�Z���0���
�>=뺽m���Ͷt|��4���]헙�<�5-��$�¡-'�y�yx|ux�[�q=�y����;[������hn���Z�����Yg��9Fm;_�OIR6Yn�����Zj'D3KptD�������)��=��
=�aE�r`t���X�"�FZ�8}"b�k�]�{�v���� )c}N�5��
��h	�=�p��1A����0��k��2�� x��a�څݥ��`K�k v�cv�(bPK�T`RlD�K�o�q��>�-�)_<���8��o�i7�T�i���C�)�ɼ��?���Na,�)ѝ%�:�-��VT�m�����y�~	R(r.����4��
�w��!��,[��K^�$�
����~�- �
�����g�'v(�mG�3}}=ݷ��J,��/�"�I]�����u7H�g�ё�'���ץd�?l+�AZ��;�?%����zsk���YUD�-Bwt?��T�V�G�$Eb璨hC��2Fh��KƱ�:�k.�o;�����l�%j��{�����u0|��"�Vw�Nފn�?�86bs��E���aa�D�i��W+άl���Q��"r�����`�	8o�$���5�e�*>�n���ݣ��>�k�qo�>�f-P�=X�1��f�U;^�
t-sp�9e��@Ժ��7#6M������$/(���3)<�̍�"'e_B�T���נ����`���*�j�Sq]\�����\}�KZ8�V2@H��:51 �օ}�*�gKڠ��V=a��4�7zI2�Dz
x4NJע�<?�b�\ƾj�x�P�G�a��BsH��X����#����PӞ�x�o�)h�@*.������
b��ʩ��Y1RY4`��<�T��vz�k�d�V�(�{�*I]��m�2mJ �r��,�����B�ad�3�Ԫ�l}}^����(�`� ����)XE�Na5;J�)F���6M���w�$w���*�͆3����r��;��t���Ca���*���JOd�H!G�I l@+�t�|�/��Z'��(H��Ӊ��)Z4�t-���j�#6NEL�;S��$~�C���UL{�2f`mq�E]S��%���9qm���U�&����+C��G��l�����vIb��!�E@�C*�-N��ڲ�_�D�Y�tb�N��Q�@Rs��(.�Xε\����'�{��
����CtAS�+Wb�f��^�4�&��-Ay�s��\�i[����eӑ�Am'�wn���v��ʎU<��L�$�A��%wQ���՗\I0-������u��S$?�-���f�j�+#�NllFvI�"�
!�F3������3d�q�4~��A� �N��'���[^�	��uj<���,K��38�,�����~�*5^��F*Ac\���sdE�ۣ�;�*"5��vE$Q�UN��yS&�nA�3��hf���v��F�[fL	nM��Z6P������f�����c�0�a�X��j�X���vύ&Mi c=g�4���}�o����Z�����I�b�Rc�{�9r[d�����U��>��#���+���D����?Yfzy��{3u���G�h ���]l1��<�jR%�m,��YT�^���"6���P7H�F���� �2}5�J���to����q�^�´k���� �ܵ9�m	c�ɯ0T�k�U���&y�㠛
xd��\1'�(��ӏ`@ e#�~�g�
\��3�|��׷o���}��A�i�O�ڝA��L3��.��ZEF�cAN� B�=�
W���Vg"��I�fBVC�p�����l�\����
V�}~����;��"�� �!�.���r�����4��3�#���5""0���DMu���D7�������
a]����S��~���H�Ň��-�h�I��������h!^�֐ֺ����3��%kД��ߊ,uk�
0=Ր6GCz�-�f�ھl��չ��\��q��=$[�dRw�eD�.��v����Xa�W���BV��#�IA���W�,��F(À�B6�׿����_��!��epTW����z���(�0� i�8�,��v���~K�K�C�)k�M��@EӚ�v��yV �JX���i�>����� ~���!n>�}I�P�.y�I��4��𢽑F�[�=�?M��.�����3<-�,�X+I/���|��-���/E�� �1"�Q>5�Z��� �y��Fo^�B��Qqvbǿ���.s��6��s�7#.Xv�4��&nt}��cC�,��������h�U6&��%�5/}g�v���rR8{8��i�+;MnZ�������NTr���|��BX�a�6�/�g���v� �Ɛʠ����_ٺ��'��0����D:w|� �5��Rɜ؍�����j�w������*��3���s��a��"�b�BB�tPp����q7v��-}��e�ޖF�U�	�n����.�F^gHm��ٮ�^���4&�DOpO�	�@}�41� ��aQ�/�R3m�/xH�lU���y���]����J�}6F�MG!ŒB0u�av�?�K�jv�6�)���ӎ�X�t�x�U_Nl��#�kP9X���<���I
iH�s�r�w��J������X9r5�?����B_�� >���S�*U#���taJ^Q��pt�SMU�bHб� 	�\ca�s�ĜGG�]��a�M�kt����v���ξ:T�</��:�-߱�[Y$'M��%�0��TN?S��I�}�O����u��1_H�P��;ּFڨ�n�������m��r��u>W�5�x�}l�G�P/�,�$d_��('���T�H�9��f�'�@�.�)�
"�1VZZ���|���L�-(J:v_���"'A�*n��% DL�f�x����vͨ�䪥��V��cG�6�H ?�%˨ɬG��z����l�i�u0�c���n�,ܒ�'r��:�}a���V1R��ƶ��e��ʀ�A�F��ΛH��˜@^\��l�0j�j�
c��T�;1�qX�+�?z��r����j��}ez=ŻP���vu=��C�����%��x��*(�	'i#L���v�Z��yQ�J�����S����eU��1W&�;�D
�4�A���K��~�0!�o��À��|YF��8	v�\��y�� ���^u9�l�1t�3���!u�p%��\�<d�f�U���.�Z2��n�6����0�L������X�t/��eSƔ48 �c�ֵi��o�o=�:��f3�$���C�<:��¢\��n�#5�w%o����$����ڨZ�,=���,�*�`�-8V@6*ԌGo}x���C1	�)_y����Q��R��@���U�� �#��\YR�z=�#	A)J�J��ǻ�i+#�"�al�HD���/�5�@������؞���|���W5$3O�YaG�@�Dٱ��������h��/n���Qg�-ރ�]��:�&r�K���$�p� k�D�R�}�G5P���{?>����5]}Ā���Sf���:�c:�>��rj"e=�n2�&ۤ��S6��.<�~"#p��q��&E(M�r'˦�5��]���g���t��
��5͇�ei��aV�j� ��Z� U������c�97� UM�{�QS���
	�Ά&Pr�?���s���ǖx=_z�kjt���>a�G��#>�u����ļaˢ�E?�C����f�&X,�RV+�l�Iq?���CF���m	+�#�����W�L ��M�R Q�6��X_�k�1p'�:号kR��dǦ�LZ�}*�ըV����i�W���i�Nၭ����yz�y�$7�Q��	N�~k��d�u<zZ&���@XK�T!I�e0[B�.*�������?�@�cM�����E�����P���ia�ڄW8m���t����v�n<�ԅ���(�'x^�h�b��%l��D���&�d���6ˋ=�u~�$~2��*�� �K Х�m���}a�����$wu�e��1���L���(ynf���> x�a��������U���P��FU���b.W��Z��x����7Q��UP?���m���Ȫ-_s`R���3_�/��ax���N�㜋��6u6�9:Ŋ�Vf�4�:���vŦ�Ё�%��00l%��e%B>#�%�'`Q )IPԍ�dhRG䋽�>~�P�:�?��O�>S��k˥�H��qp\8`l{��-�.�NV!f�/��j���i̲*���!>.ݕqj"	w����K^�
t�̢����BK=� 5�EPz�\���8�̶�P�����7ڰ��r��x����#*��öݶ���m�%vT���{���UP�Ou�A8a�B����Ċ�f��C�HAc;(���)��)�5y'����S�<�'���6t�M Q!z��ff�J�2/8���t�5h��Y·��04.��HW%�_Z_{EeX
� Ɔ�C�o�T2�_���&���A�H}x��'rN��pX���.��}}yj.�0�k?p�%e�^D-is_��4%�K`�n����D}�M����>ـ�s�UQ�\}g0�����*��&+e.e�X�X�F2���ɲ:N��UQNbm�r�c{$8�4�R�^~%~Z' -o�b0�q���x�����&ܟ���WU[t��Zc�=qWR@��w�:3�?��s��W����g��F�`S�,���sI��G�M�	HZ���_�ϒ�"�Z�9�3�<޲ͻ.� _�<c8bj_dШ������E���A���r�.9��"�;���+��91��yq"����4�8�����b�B�=jW  U29�Y�^/�l�zȺݷpX1T�x~��C���{�0k�^�fG~ 3>.��?���eq�@ ^�.�	�n���iA^}����+3aa~4D��u�W�]�dC�\:����\�q*X�=��0���E<����0v�y`V��Ҵ�9��J�ȫ6�p� ��M.�	V����g@�����S!�L�"�`�uS�pՓ�i���Y���5�GY�H�{t�3c��2�(e��{.L���~��;6���sC�x��
f�.&���D�
�ح���I��7�tg�i�[�p�����D$dB��#1/����y��3��%�ڻQqF#��ېᑦ��vs&�8������!Z��d��ԍ�J���j�=�������h79I�}*��֍�ЂԾ�W���LUwE��.�B,V���e����7c a��wI���U��ս?��DJD��@�Q%�������ߓ`��&FyAU)�r�6��<��xT�@�ׂ�0py���b�5d#��[I�����n�h��	,����f�1�6II���#���8���a�e�2w�����ש�ˇ�z!�-���I
fun�6a:�O̓QՍh%@`�o�tsS�%Gsk�cHө{��8�)$��f5��x�����s�ö�ph�J<�g���T��C�<�:�>���
��h

��������&M}�m�=�� /���X����@|��cah�j��a�ŶH��ꪙ�w�Bs-�~$ܻ&(�b{���0d�����Tjd(S�e��[�S��e�C��� Ġ�6�����Th&(O@?vrC@	�7�<_\���C�WY�
�=>��&b������6��gN�6��d+E��(�D�iK�h9ت*�R!����j�|#��6�d���J���U�	����Wb/����A��B=��,EY�_h�¿�&;g��E�@mz�VMRcQU�h�x�$�Q9�5dԠ���,����U#n�Lb�:���*5 �� mo}�e�\q��a�r�K�j$���+}��������-��[.��o@�����m��Aݝ�ɵ������ayl�∗�D
����LC�W�!8e��uq�r�(W>���j�>X�#�w���Tq^{@�4U�W4DxƝ[y��90��@ʮW>�Ӻv�ۈ��h]�El�X�%�8���sX<I>ї�z�HD����AE�䮒ڦ�z�"+e�U�ErC�,H*%FB
�C<���=͜���׷�k�냺�F_��c������em��w�<wN�.B[F���� ��Ş"�q�<0�|����D�/�u-~W�2i���Ojk-P=�f�r�=К���F��na���^���-�#��}��v6������G
Q ��{�q�Xm�P�dlJ��)�}�z��@3�^�܄���
���/���z&�
eՕ��u���i�~�0�=n��k��+������Ƭp�>��C�t�E��ǎ��٭�fH'��S<B�l��h�B8��'>s����yC����A��}���l�=.�-ܖ0�)��B��2(V����Q�C��f8?��m%�/��? ��[:X��y������(�z��8^�s����=�P55D�g�Jg���s�TC�Lш�f@bYY�D���$ SB�c��d�c;s��m����k��b�t��Bg�,���n��zn���5�K?�ˮ�oڇ�F������A3�����d�Z�u}s*�_D�p�*��8����E뜬��ؓ&f8#�ޒB�xu���g�$����[�ƼYrl���:Q�vO)W����N��l�@v
	�:'
5��Ս�ڦ�hр���c����Cx�� J�6n����u�4:��ƴsе��j�h��5#ѷS��ᓧ�<(ވ����k��X��k�'*��M>���r�n��x���b
�@Cpt��L�LJ�����#��^f�mMY��֍{5��P�4m��3�$k_H�_�T�.�З
t�U�ˇı�%~�̛ ����� B�3Cp��N����<���(����VL�Ҡ�N�r}~�R�.�O�p� �������|+�(n�=͞ǽ���79��]&n`�껥]��$���%��\��U��<r�!n,�L��wgD%R�Jc�y����W�����hԏv��q���8
���@#��/��^��\[��Y���\̗������jh�ۄt�n$Q�'��L��j6қJ�/�&�o͖���X��1쮮���:썙Y�������� s{%����.g��Ò����Pu�|�w�c*�%K�BԘ��&}D�o</��ƞ���|`������ύ�2��yKҝȰ��
]S��T-�����ӏ�ɹ��q�8.ǇB?3��=<��t�64H�\�s�j��D�n1�t��gK��۵�X�`O���Z� 5�t�0=ө�M4r,�)���<.U�W-�L�K�k��ǯ���Eo{���׳��\'=�i�W@dd��{��\l³����e&��`�˺�R$i'�q�,@;�r\�i�}Z�H�t�si�ed�a��I�}��/-i�vmrJu�y����4ბ���4�ME��꯾m�3Tp�|
�I�~��]��-a��Y��o�ϱC�G:�ߥ�q���g�0 �f���_%�%�-�V�XJ��E��MCzڱ��D̗�)�^a�m��0�������C�=��->��1�.�m�)Lيͅ?��D7rdc7��oq٢N6�kA�"1(5[�?!Ĕ���wv���Txc�y؜O`���g(�ѹ\ȊP��F��G7��^�[���ů�{E�%�
�sz�F�������4YJ�𛘇	-Z-��t9E_�j��ٕv�uyz����/ȹXd�:$���z}/�q;�<�9��:�S�[bjZJ���p��N���)���8���k-@ oB<�0.-hS����_���n"խ������j,k�:9��.{��%DJ�F�B�/��M�2v�D�E�)��J���Q���O׿����Uƕ!����>)A��ژh #�mcA�Y���u=�$�F�^d�Ձ)k!�2�j�>x��Ty�˹(UG����K��k��b����f;�z��>3gݵ����i���]1��Q��d~�c��ZUy�O"m�s�����^l)����xU�j��Ey��/_b:�.H�Ll!������oOq�BJ~�����W)���ڲ�9�`:Ԛ�f��ᦈC|���R��鸂,�g�~B�S��T�v��������Bl9�k/ߤ;�[�a|����3w��-1 9�hY��I����`3J�'sRx��K�a����M�|�������l�N����&��py��E�r��K
L~���2�^w��xi�wA�*6���d�[��_6Jpd�)��i?�H;����!�S%cQ���DBU�����C����'���H4�бi׋�]s���"z��Q��*�v�&/���Ч��3O�} ��z�#~Ky���>.̤�%�����!Eڻ[�P�y@��] ��~�-�b�Y��\�oz�7�f9�֬x)B��؆�����=SU�iV�^�,ϱ�
3�?�fJ��mD�%<��|���
�L*=nwh���U�)��L�[�����k���_Ǜ/*dk.?JC8E�!˒Ƌ��E�d�_Ъ�	�c^�	��댰�P0TR?��FW�Y�)1<BEWM��=Z� "%��t���b\��D��B��b֦V��ԕ��O���~�2q`�su���������	 V��X�G�c�_;TҥcYus�eJȺ�Or�#���2�r�n��\C]&���)�.��ys)*Fܵ��p#�$�f��(�8�s�5�ϖ���<������z�R}�F������B������'p�����F_i��F��NT5_�2/���}������������3�҉�y�-Ʒ�п;U$k:��1��_+�`�-�������_�E��G�wt������\�;�0_�#B��Γ�&*4Qcl�i�����g�#�WIݻu^�
�1��tܠ�uXWvI"\/v�K)�3W��Y��o��2W#m�g��9vUeO�h��,-�x̴}5s�����X�%lŉ������#o�7����>� �J�FͥQ��g�x����tϞw#?<K@�ձ���v���]�������NHtt�f<�(P�Z�oi��$�7�^���!��>4�N\V����A/(n�g�?����c�$�����+��ơn�0\��e%89j�Q��(-j&��%���Yy�����͛�1�S*I��*2bN��@q��R����B�]�{hy`��B(	-\} {^�.:��6c�g���D�ư�'>�H.�=�s�h<���zp������5�w�B�q����`�Ʀ$uۛ���yY�������Q�Z.K]O������)�'�vB�7
~��m3),�P51�ĉ�Q�Q���|�ܹvӠ(��!B�y�S�ἃ�9�+z���N|H���S�q��wN�7� �ÑZ-6�$G?�v�ŕ���B+rr��;u%h{}���u3�P�8��&����P��9]�2g� ����*&�L�r�{��DL}g�,�0���#临�n�2	3ap��BZ�v\n��g_Ƈ{#��ԭ}�u�<o��{b�r���RϢ��0��v F+0-�'�v��дq���)y���Wϗ4�25&��<��T�Y)M�+�'�F�:�>���3�?~�U��Z�WhA7���te�����?x��CI�D6��MU�(w�c�yT����|�n"E���a�a��#�y���L׳���4��Bj+��wS�5��������A�m	Ł�Vc��F�=D�x��{��[	} ��-�_����)�L*�\eK�e�1���ހI��M���Tco���+K���"|�Y�nZ��Z[F4
��k�B΅۠�*���-��0��ݸs���!u�f�Ij��C�/۷�A�(,,f1۹ڄ�'z	r#c8��Z�-������D�L���<�!
��3�r)B��(�%[[.9��I�m���r��8}��6{���rK�u�B���;�LX(�A3)�&�����d��S��BF%��y�#�D�>)�W�<�����Սx$���a�Qe��!��?B"b���E������& J�a�?��/�`M<�e�>1��ŧ��ub�d6��<zѥ�+^�j �W�����1�M=�C�����+=eY�)7-l��8:k��w���f^�N�L��9�u]9�&]�yk�_����^��KNB��r
8�9_m̻��;�L��x���%iU.�<O���:���m���~)�}?���s�F�q�͔	��cik*��O����X
KR͜>�d%ІA��H��0�`-Y��cl��WE�!�����s\�q���4�*��o�
�R��#k1�LO�����i��3\�~U���K�3�]����!怿��͑����Cb���s�zy0��Ԃ�|�E����$#>��	2�]��.*	�s���b���L��8Ex*������k�'D �b����+Y?nq��&���x�gEW��;�/�=Jħ�M�+�G��'��܉��MJ;1�{�(Ka=��U��x9-w�׈�*f,�}�Z��?�j��7�5w/¨��	Y��G7�c%~<,���A�;��|��{����\U}5PQ��
>0�(sǅP�g � �l����_?�` �@Kb�{\#��_�y��Y����'r���o��W]t���0N�'�g%���J�Jʅf�j���B���\���)�{�3mw��z�P�+o+L1��+�e3e�
�s ��Yà�hN<�!�8�*jP�Y��A	�$�9��\%x���41��gThi�13+l���AH���-���[�`�����j2�н�?� :t�?n��5�)�
P�FpaqHR�+O��)�8Y�7��Hɽ�Z�"Y�.9=��l�:�4��y�ٽ/?F#�T��t9Jp�!�3���RA^�h[,B��+�n�|a�Q��f��&l=� .�G���p�7y�[W��L������a&�Pk�B�񕱷õ%f��s n�o��P��^�W�΃����Ա~�%H�c�/*��ol�O��3���+��	u�M`%�����	۩���,�%5�H#.v�3�[�Qi䳡���a�1��0��	
��U�G�E]�a�,&%<���)����1qJ�&�c�'r�@2����.h��)����p�0�EL:��_�4�`{�ڈYGx�7�w�zHԝl�|�6�B��1A&�k֙`�	sr�g5͒ư�	������aG:�?[T=�חQ�6f� P�M@�h�Q��f~q�%w4O�0��.�w�
�����%��M��-��V�KO�����?��\�@K�������Sn{��r���m�sU�A��s���E2O�U>�Y�sxLр$�-����+�O��]\%<�,��j�ǌ��QO?f�(+�ko*�{�C�dC�,A��U䩲�@���� �z�� �1�=f�=�m�r��՗k�N �5�_XC¢�'�;���4.6�5&#/r<+q�F��� �7��E��0�r���M�~���ƈw�\51�kN��m��N[��n��+�$�d �7�3�&��A���&�N�\[ �N�39�]U��{�N�ԂXgd���������R5�Q���0p��?�lc�:e�r����c*�����$S�̆���7�̰��y�ɨ.I����e~9��F��1�?�J���T��ӘсWf��8�5hu��)(ڜ���1�i�s�RPiӘ���|�!��hf���]�\�v��a�b`��98�ܤ�.K�a;�(���P��K@��qIq�!,)�M�Kcmy~�Q�%̵�	�K��c~�a�b]��ڏT�~��I3�B���wn�	�p��O"�h��_㺧�X�M�7�T���j �Q�����^`���B�Y��^��fE�|2X?q@a�p�>֯CD%(�W���<+c�U1f%�8Ө7=�#}FYi=`8o�&MU56��z�6��$@ܳ���渞��X�h��)�3�0�5�2ۉ��D(�"�59ׂm%��uϝE�E���% xNd�E_^�1�2S¿��HK�?t��7�	f����-ɸL��#@ck���?�w�H�<�H�{�/	���q�4w���bM�:�r-?A��[
 K�e�=�����F�@�F�4ҋ�'TXx���kV�^�������&��'$oY�H�,�q>�D6$��b~P�"�A���EST)�2���؉{���I��wbߞW��9/ _3�7�|#[�FV�� /ݬ��Y2�c�ι�[�'l�׶+M�+���ҽ��H{����Y^ �߮/�G���pۀ� ����+�#(��ZKE�P��A7�r=<�jN1T���A�Y�PZ���_�4���K6��FH���8(�	�M[�{�htY���(�x1 M�D� F�$��9�ᘁԼ�|��^�h��
Jϑ��w�15��rl��_}l�������'��~�;�Z�h���c\,	}�E5�'՛B{l�E	�^��k�' �l�i��c�=h�"4�A���o��W�%�\ة}��K��f�� �[���|5ok���_��^]�n88���,�Sx��"m�����!���u5
Kю���z�����FК����ߝ�)c���Y$���V�֒�u�k5��nbݐD��Tt���Z;����B��#�DS�R^�Y�NK'ԲX]@�8l//4�dK�=6!u�]gř��wu>�=�e�Q1Rx
��4h��鷄�DN�Ok�?yG�9g�;�r�PcbQ���+�#������7��h������O�s�'>�p����:+�V}���s��倆�����W\��m��#4�J6oT�}���Kا	$.'�q�_B�N�A�	�V�ܣ�Q�#�y������Zu��B�x��X ���̈́N �{R��s�C��;w��r�����u�k�P�f�eh���?a����c}�{ �\a0�Կ��.��	Ƌ�D2�F�$���W��@���qʊ����
��:ƣ\�2���m��	��c*2�]
T� [�U{[���#I��cዌF ��ŉy�r���2^�y�v ҄A%COf�0;rUR)�xs��s+_�jh
��ɓ�]�B���_�"~Jj���;��'���R��`G˦P9~C���t��㺛k(��a7=�#ؗY��F��L�g�%�'K�;�y A��DAMc%'�^��������p��Hm�-�_084�k�~F$E[^ 첨 I�*a'������ջ�ËC�H��*���X�n����C��W��4`��3���F�C���C|[��� �D5��RV�!�aX^�ˡ��	��`3T�~ܢ��`i|F,!���=/�A��m��93�3.�1��z��?��-{�?s-���k8wJe���igv�O��\�����^R��A��I�R��U�"2��>Sx@"T<����v�bD���}��wAo�,0O�'Ζ̔�� nރ�t�Α-H��Zр#�=ܖ7e@x�,K��
ӳ����,����>h>	<ǮKʆ(��k�tN���GЈ��	���T��T{g����~A_��5��5�$wyZI���H�cW�گӲ�qo}+��&��X�s��kX�2.���ώ���9���� E`�����n(��e%�6 ���f���,����"�/�Y� �=:��F�VϚz|�s��Q5y2���Ak|���	���"�A�b�5:�u���J�7aV˫��3y�B㾴˨��Ι�%��&��	��e���c���K�*>��"}�j��re���gx���%3;B!�f�s0���M�n\z��pع?rT�af���t� h�25S,y�<h�z?o���^��C��]�a&������h.�>�#D�s9/��?1�,��e����B:bz�WO���g����A��fH��R�>a)����?��i�)۝Qĉ#v.��Ld���d�>�����ߕ���������ٚKVr��5I��f~_1-��/��ź-`��z�����h*�v���)�o���#d��'brv�yR�A�V���܊'2�cw���m�7,�Ec�H�^.b̉���x,$ȝ��{�u��6�Hj7�b��8�'`�'��w��.�����X�6|�-ݚ�D��3�t�|�e:,'hdx$�I�\Kp��'z'���ZOC2<�p�+䐾�zXR������#H���Dv@�/�K&��3��G�*��SQps��Jj��� �:��\���<��Aq�W��c)�|�6a��F���B��	�9����/�}~)�2Q�I$��?��eZQ7^�;��^��F��H|��`�^J8e1x�wq�I`M1��������.RNk����t�)bͼa��������Զ���,�?jȭ|�#���З:�z�������8����(~s<�&��@��ī&Df(3�m��*W2�sU��NM�c �ϋ\)e�5�3C�)ƥ�^'��E�Uˀ|���K^�d������2����F4��^a��+��J��6�L���@�g\n�y��p����?�����:�UT�x�]��9��9=/���s��p���x���V���}��1��A����3o��)A}r��	�`j��"?[�l�)��/QJ� �Zq�v�_?O��v
���#�ωNÀ�.S�@������^;ĳěB��ؙ5J�T������qxZ�U�~�x�Z�(ހ����q��¨h��Bu})f����e�Z��dN���A�>Kt�Tg����v�g�..��%+�蝖�}��<�9�q�C0�N))m�0�v� '��TA��^e�`y>�up�K�eD7�"�JP�>M/�,��b
yұߍ����'h+$�r�d}G��W,u�̟�)_Y�\��B������&]r����	HR�Q��Lؘ�������.1'à���ҫ-��2��r���`�)*i5��JN�Ȃ��ϊ��+c�ނ��s�����d���`K�����k���I���X-P���R��0� j3DJ��=~��$^����;?j�}{�ŗBX�W�\�Jn�� 'V�������>D�=ͦ������ǧM���^�h!�NE>i�+��
��ojalj�}s�ǵ��DEVu��uJ��5�ddwz괘_d$�DR�:c�]I��XDeK�?�˪c; f�kh�g&.�iO�~�[`5U,{Ţ̒����M:R���L��;KCH*v���N6����kf�j�Գ��#~2ܑO.6����غ#�i�����z�lgݺ�M䚓1�B��so� ��?Qp��cz��F�S�K�%_��Z�G��ʻ�+&�=�\��P�gZ��0�.D��΍���
�C'���M��[bAc����@5�G�%��P��$O��?h��T�Ĝq��e�Z��@y
>��QQ�i}w��T�<�9���#;�<�!S���"��׉�X�g�=&�K��'.�s�@��ܩ��g���rHf�d��q���C �e5<3:�D������C����_��f��P��S��5
M�JP1�Ċow����麌M�HIhp�<j�[G8��(!���h�[�4�,��`��qS�V�"C;y4�������kw��H��N$�5 ���p�7GU*����n_Z<t}�9ss�����Az9�4wIw��k�aD��K6|1���pɍR nf�yn�&Via+��U���^̸��N�H�����Q /RU�0��ar�#=	 �(�e�E��D	����`�B,9�h��W �p��G�'T��1���W5D��ٍ����r�L[x��+����o��4?pL?Cb�{�	�WĻ@��`�p�@t��V��8=��m�7�^�0��8�ݨ#� ���ڳ�M�]|2�L7�Ø�[���E��g���7\�����AHȀ_�}(�Y�+�S�~��g�=#_ 9�j壳jP>^������8�ˌ����U�����n�+0�=ҢS-jC���?�Ƈ�zN��}c{u|�O8z��������aZv�DW�>�Q��Pt.�q$��g�;�����48o�O��;��uF����&K���9��(�4FI)���$����w�]�ǡ����Ĳ�n>U�-�������D�+�W��Bqϯg*N�I�<��e��kM� ���6�DN�6R�F{��P�@	�<�&�ۿ����ˁ����Z�b��=V�,!��]�~��R��eO��b=��q����Xa��B'��re ���Ӝ4~)+��\�!�\�Ĵ/).X@`���Y?Qh���L��a �B�в�%HF9�հf��F\Z�*"#�h4^�&f��EZ� ��'_���'�rܰ��|�d�[xUu���lpV&?)E���w~���������V�mVYӱx��M�~���֩¦�s��o�id�s3��C���F��M��.���n����]���};Pd�=@�L���]j//κݷsF����2ܞ4��`��u���Ã���Be�@�����N��Иk�j�(U���zur�5�{�;�p�fT�rXL���)?�E��o��F�j�W�Ŧ��\Ρ��q7�jy�Θvj���B���ݒ�L�=��B�Lf�0���� ���FJ�A܍2ٙ3L�f�)�ӟ�m���7�$��>�k}��ғJ���ٰ�*ų�Vtx��,����b�}O���B{C����Kd`��p����P���^��C[�T��wR(>��^:m�����Y�@���֯uםSC�Up�hݸ�LI�O��������^�aP!Ya���2���~Jo���?!��I�2�®��*��8?��4�H�Z�L�	����ră�"U���"�b��7B� �J'i�����7V2�јKW�b�ГUK��4d)�����;�q�pYXd���ާ�)�`yB��WĮ��~#x���D��$�
�٤>#f�W������������?�F1RGa�66-=GV��0lB�P�BRB������ty5k��n�z���1��]G�v��t�S;L��&�s�g۔�Ŷ$��{f�p�"57�7��y�����s�c>r�/����c��X�O8�ӜVP!A��+褵km���w�`@`��zb�3Z%��e����!����f�p�kYrp���h{��̯������Wq��U�xN��_�Vc�����M��Z�|��=���6^h��{$ �jz���3,ؑ,E���")�*��ى8jg�Շ�c�װRd��y���)8a�)��y�QX��t�-�$�ջ$eԞoՕ�K�t-��W�2�vu)��DKJ�F�o3Z�0�銥�ѱw7�S ����!�o�q�F�6�q��ͷ~�BڮG����J{�z����
(��N��Bok����f8�)����w�$9H"^*)0^�;�'��Ҟ��r�FB�Fa�]�K�թ�/����埂o!�&[,r=�B���@�!A5y����x�ۮy���у�u�i-*�P��Y�]]Y��]�R:���h��}�A����$��i���栞G�۞�t�}pJf����?�\IAԞ��QnʴΫ�cX�}��wd��(��8V��SOA����f\�.e|�x����3$�$�U������u���ҠP����M�� �*c�{@/D�^MQ:B���t��H�z��pF�n)f�߃�<=���H��_P�@����(�� kU���A�Qh�]o�bfoߣ��k�EO���n\����]y��Y�Wx�Mcgpm2ۓ�Jib*���hMND�Ŋ)7��������Ǐ��x�1 ��Pt=��8h�Z���� �0t:WO�)%���°�	�]�&�¤�\F3�����H�����\d6�8���gC�5�a�u�8�`�B"�3��}�G>���[c�=�ݬk���\Xy�fko]l0F�H�c��,H5�RL��A>��~�v�EF��M;r�/d�VY�k��|+�h��&�V<&f1�&!���7a�R��&��$����L��iݝ7��U@��C�	 o�O����1��8І�Ӕy��A���>-73I���v�߱�F�ֱ!���޴�(�/|�7���8�*LS�� �K�z��I3�Ҧ\4�]s���(TS�<O��DU)w@�8�����N̔�mC����A4S�5ϵ���dAs3�c�յ����� ��-�r䱵g���^s8�=��D��cgz
\�hh�I��w�u�{5R�<�8��v,R`���b��od݋Q\�.Z��Uwz�_B�1\�d׮�&�����3��uz�mם�2���n�'w%ج��U�!z1<�l?� ��F�O4����ڏ1�"���Q���d��'�P�Z���0���"���(d7�yn�Hs֮���v;.��2��&���
e~0<�� V#�D`5^5Oy_Hie��g�H_������:��Ȏg�]h%~�tW\��B��o��t�5 [�^i�>뻾c�'w��\���vЕ�*�����b�tt�w �ۙm�fk�w1�4���%��x��7���Vx҉^�A�fM�?��5Li!�rb6��ID�7�!��8Bk;<;�4
����}�S���M��E~�!����o���B�N�+(��G?�z�L:7��~CG�\�}t�X�k�F��F��LN�^�����W�g�"��_d;9(<��<�3�Enf��߰�k�1]M;��wM �	�+/���d���#��`��ϲ��}2�M�Fb\�j�����G �9U��	��e���S�9&�^�M*3��8�������卄T���y��7����0�^�,�����4��f �)�e��p_Cik��5�\��8Ѻ�_@�����m��C�� 욪2L�V��z�D2��O4`��C8.+Z��91-�U��v�r�t����a��K���x�*�VN��*�"m�
�JCUs�h����Cv����D�Gu�d1[,"�*aK����7�"@B}�J�D=�1(��r����ScN���$|+�Q�'�sжy�g�=�=�����<7c��l��X�6���uD��*F�#�R���VU�\ʖ�m6�yP��A0.�4z�NH��}
��o�6�E�����C�25��"���e���&d�;�ݳp������,�<x�$RX�%D$���O���wYu`1�N��V��ڒ�)q�ޜ˛G����~��G߽S]�ᒞ�  es;bx�R��k��Z[�����=Zx�_1�9�Y Z<�.�W<��A{
�6�oA�y��gzL����c-hn�಻��CH�9���ws����ʛ��ǚP�84����.�J�2Ǆ��|�A�iG��c�6�tky��*"Z
�Ѡ���x�8[,��}C�ȯ���A$�>L8	��/ʰ�Qʓ��מ�<����3F�ݐ�B1��' ��z�ϩ�!2�Xn�e =5{:N��x5�,`��?G�D����P'b�����+Rĺ��?�.΄��eN�"S?��x���|[6�Q�,kТ�w �sH\�U�}�����"�.��Q� �p������Z{�/�3�0�f���M�<�gg+Kx���Gɞ�ߟ�/�x��ߝ�F`�l���O�Q�fR�q�㗊����$J���	{���0"`��sc= ��~����J]���)p*5k���O�C45n�٭�������x���S6d9���M���pmEΘ�H�76��LD	�}�b����o\�Ś�wq���%$	�{�������@�B�A�e࣭�<�!|�`�.o>N�u �ٓ�f�a�Dj分,i'�ii�
kr�KH�|���΅��G(>j�:䎅�;���BK��~�Vǽ�dg�+��z��E��qg�:A��h�֮�Ģ�#�9KZ�m*Du�����:�N�M�v�0��y����E�0�Xv4�ya����0ބ �@P�H؟+�	2��*�a&$�˶����G슂��͔��Ь��ٚ��s�e�Ǜ}\��F�i�Ͱ-�@��N̺	�_�U����<�/ԏ��aŉ�ZfV1�]�_�0�8`n���S�)�����'֘�Շ`w���M�pEA�ʤX|��+ ��A8a�© d��i (aŴz\���$���*����R���,��d`M���a�� ��T�_9u,8`���G�Hx+�����C$
\�g Z"@DfO���ǅ�B셠��99mi\`dpN��g���c M��8�$�^��$�2�&��"vI&��R>c4��;�.���VAh��1�vT%���]+=��Hn�����{�e��2 �����B[,�d�k�a��ΊOe�b�tq�C/qn��>9%Z̓�P"a����w$�$3,���l"�WNI։��Tȥ�J`�SڎW9jY�g���9?&���n�4�i�o<�o�ƪZF##�wq���f7� �sV�B��V��_��Q
% �ى���= �ؾ�]�	�jR�ȡ��[8k�@.2�.~z���ىGE�� �*p����� ���/P�t�e�mؗ�>	��dtj��˒�n.9~�.��uk�,��ڌg�{�&�(յ`�{1��ƸI�-#0��[�*ӄf*˅��ڙ�(�F5�,��ȿ�#�<�@)Yl�7�F��'����H�s~�30��f�uJ�W�2� }XΞ�?C"2O ;���kV����Qq���/���dsk;�[�Ǳ�H�-vx aO*nm���h��՛f]DgH�FVޔӫ�p��p9�XOQ]�=W6�׈Y���<1$���5�.|����#p�q�/y<T����,\i���}��B3�����l5Mӏ��7q@gb�M�ذ��8-�u�a�đ�)An�1ĉ���w�X�����&Ut�f;!ڰ�'�yBP��� ��9������}{>zI�HG�럳���f��ӋLӌ���>��r�`e�2=D�GU�Ju��-ʷ�@~iȯ�dn����8C���a�X<�P��Ԩx�%�_��0i��������i�df�o=:4ʾR��1O��@CPM�<c*v�E��EÝfB|$GBHr!wk8�u|�Kͫ�粿��).yr�}��� _����[�*�ie�@yp�#p���A��\�q\�|�~��%*�Cs5���� ��B+�fݝ�d�9�}X��9�D|b�WR�����E�$.U׏�/~�6�|m�����s��k���T�̊5uq>b*�3��B舊��<gσ@F�<�:��eS�[4���|�����-t��_{5�����m����(.�a%�I���E�7��gE_Z4}�����l�6��pO5��X�I�y�9��*�7k�:�uBֺ�E�~Q�ڌ1��y���5'u��&�4����B�Q�_����V�-sl��ް�V�>� ��B�  q��o���CC�G�;'cUu~�ƻi4ZC���>5��W��kb���z��#�||��\�-������6�
ܦt���?���ġu�#+]���gAm��s��5Y�,]8���8��4P���r�\�k�  ��|�&6)��j���e�j�i��c-A�c��#��h[tqo�(�>�t���Z�uM�j�6g�+r���2O����8��	DĬ���'u�J)[�C��;'cf�
C��pZ�Q98�Hۓ���r���D
7��K��W7eT�2�d�$����[�öd\��:��d��h��7b!U�!��F�7�Rǫ��jCD��?]��;�`���<�ùv� T��T0_� ���Y��Py�OqK#q�~b�y�n.��'9���2" G��X�)����ػd�����29I�4=�-DVP��������_�_�S�}Ov7ƥ#K�e�Ǯ(:�R����$����-��-k�|F\F�3Ia�^�U�Gǥ�'iܸ8�[p^X��p��d���
����K���۫阡�i{��'г����sH����̈�r�H6)�0�c��M��[0M�`���Zۂ�k�������_�?{�K�W���l���%�t�/���G!�my�"uk+�<w#�8������އ�X�(0mgl�
 �R':��x�|����{A���4�w�4n����d�� �C�f;�`�%yJ`�'��$zHh|o��FOU�ڎeA&����΢��Γ��\�`{�����k��Gw�Oa�ew�_I��:��9D�[+��s�^�
�{N���Ab`�t��;91<g0��y{���RE��73;�������v@r��_�z�0���מ�L�M�C����@��okQcL]	�4TD*8�G�mI�1]f��)5��
kl�'{x���6r�������vy���Z�	<����7\jVߴn�`$J�G:��j&qW!�j^����yd�Ɏ�:;:!_ո�9�mҥ�i�s�~��o�����\~{���G&S\��{�&�[)<�"A"�I:Ӧ7�9� ���K�)�d�C�b�:�N��\�R�h���E��)�VQi�W/��30*�ڧ�my�Bt3O�oшɻ��a��ŝ�8("ʼs�)ٶ�jl���nc�ܡ�I5��+~�B�E6�g��&�i��&0̗�0���7+�Z���6����W�C��V��"/��v�Iݷ��(��Խ���{{B��u�WޝX��럈k,0��XD)^;d��As�z�Ȇ׍Mۚ�5r��=X}�66d���*:}�zX��P�M.Fu�o,|,c#5"��Z��j��z��@���&ѣ[���}q� ��L�� �<�Y��/ەm��dѱ0����i�-�b��պ{������t��П8԰���D�t�ߋ0�m���!�0�upU��Y׏�"i��ɇp�[e���ya{i ��n�x�ޚ�'!ѺsAB�Lp�:��#}}iS��	��㋐h������)����V%���f�tfU�x�*Qd1a����3�3u�O�@P�1K.7����QnM}(�r<�+A��o'2z��}z:����;��3����ű�9C�����)i�Ŏ�H�TDo*������n���\��Ō;O"ʊmf.���>B	u�V�=���]�b�fЉ��N�n�wT���#Z%l��w��{�o�ޞP򴪚��(X���Ǎdm��i@�@����1=�klZ�\��:��,=�5�zn���e�g��dK٣��Tc�z�  �l&zT����u�)�ཫ)��Z��O�R�mXT�/kI�㹔O�WGi]�~Zz��v�����G������`ڱfd� ֦�4K!���E�#�8�)��[��1�M���/��r��c�H.1��ĕi�kK�+wT/��eB���{&E ]B���$�A����qG�q#$����!a4k��b�v@^�S���[#¼��^=Q��d,5��2=h�Y�(1��T�Yx\f��Et+�� {5�q?F�]���|���:���5�h?�����L0�~���m�H����	��_A��^��l�i��7���|{�R,Q0p�'e�`�w]c�EUGdh��O����C9���<��R����v�:�i~����@��ڴK�#�3p�[�?����.��f�9ј�U�F�q,Z��e�4U|>/�ል�˧՘��Q(Y�O N����hfvd�A�}d����Λ���M�e��P΃oK�=)P%N�jP��Q3q�%���M�чG}K6��1��I�`�,4�Rw��N�.���׀h?.zNJ�.��|J���-sIU���5ؤ��N�&����YZ���#� %IL�5�XM��K|�X���C��ڝ'����#��,�N���'fWd�b��w�rBN�¾���t��\�ӶV�_~7�:]P�P�x�C-�X�c��V�����FMES�X~�P�y����1���g�S��u���'nʇ�%&����1E�0�	��{���m�����癄L�����4j �܆zL���bםS�㯲�Jp8��cƷ#����fͻ��%l���F��Oz�MxD��Fg�FQZ��u�B�T���=�p�N��"SV��	�\�Q��!��eG�z*0��8�
SEN͆?��4o�ڧ��ъ5Y���wG��T8���u�k��!͝��d��:�e� b�ݍ�Յ��L\h��GDR�/^2>���+���#6�Aɩ@��U��
��\�}ep�bC]*�l)P�y�bzjĦ�a��Rѻ�ߒ�<�'��� +��������"Mq�T��&2�@֋�)����X���Z�1Ó�H�k�$7p�q�+�>4ؿ�ء�j�,�ޏ@k�*7k��j>�an�ٳ&$�޷�'y�������FUD��� ��T?lй���PD�
]WrI]J�=�xYn��h��k\b/2C�ڣ��C�=Q�'���I�ܚ��S*Xp/� �JU9t�*��S �L<��Xd�K���Յ 0+X��l��8�.�d'�ٹ=�g���Ɠ拋������i$�v��ҟ��Y+a�o���*�����u�dS8H�6�hkA��V���I0����f�ihr?���>U}�DA5z�bY�!	� ���ӰC����ZJ�T�8�-DeZy��,-��l�'ξ����;�ҏ��@`�כ���NQ��>"Z!��L�fI=C���bZ�qԶ6`�AX9]K�;�G��_>!�C����KŠ�^8�JfFO�[�/]���p�
�CV��~/��&�/��u>�T��|o��T"aV����+�vΝ�h*�������4ճ����	���}�W�&�:^mq���P䮧��+�#�N�a޽+bX����)�*;�]���i]�Q��=JiE��UK��r��������=���c�j��EJA�n� $G�<PK��^�_Nl5\�B�y����eP%�^5�_p���$�8�:�Ǚ����U�a/]�<�A�1��A8�L��I����9Cŗn���'�>N�Ø��S�q��=9��.�Z��A�>.hIsdl�J��'V�O�=|2h�$E/!M>�����h\�P��}.��j�'�-X{)ۇ�@��oھˬ�����I6 ��� o5s4��*�p��~���d���.�,ƫ�<T���p�BZ*�4OqX�s	5K��_G��:Xrb\<�F�']���ryX ��x��P�#�K�%V��U9+���V��7�h�.-��r�h(��VY��PU����?�����&
�{�̩1�p�!��OB��><\6�Z��' ,vf���r�'��(O��u͘ �>�ʹ�dEp8�δ�H�\ײ9i�xAc^\���^��p�.�@�u§���B��P������M�٦XYb!xP��f��O��p�+���N���{����--���.��C��	ۿ-�W���p(�W���Ӂ�dso���|���&ӏ�g�ٌ�?M���P(	 u�� 8�KnZj�d k1�|�c,ϙ��9�>A�L�W���S}� :g!�{ș<�؋�^N\�`n�?%Q8�f��mi��g3*Ͼ��Q�H�,��p?[8�zW^�(���������_7:�H���W
�����遳r�w��h�<m�l���I48�܉4���D�Q�˓��Y�GO ��(��n"���om��k��ۓ%Cg��F����ٰ�3�Զ�8���+Z1P,���46����"?~�_�T0�+��V�\"t�΋��[i[/38d�=��A)lwI!m�g��ٗ�αN;�tC�ٌ4_���l��[����L������ ��s,�am{+����*���	�*,���O����'%y�!,��$?��Ź���	D�/f��[��}�����۹�pֵ�Hh�m{���H~K�X��@�B���?{r�z>��{-[��f��/���^sn��*aO���:��w��G?=?ۊ�� q12���&%}g���*z��M�_כG���EHp��8*=<�mH�g^�,˻%�(49�c0���j�����u%J}�lvFJ��%�v�6x�`��q-*Io���b�G���E0/�<�[`�����X�����K�@r�9^����6��8Ż�ג�C�Ȯʌk@s�����ȅ�"�H�bA�{�:�f��
�ob���H���Qp_ߐ����vJU࿵(�j��>]%��_�x���	�vK���"��w@�b-�W�gN�Ox��GT���ӕT�$7�}az��C���`�T9���(��)Sy��|���ɰ���'4�&�AL�vSr�s"M[{�V���'��hA�Խ�6&d��9��)��'R��p�I��H�Ld�Ԟ�R3�!M~����C�t�C1�U�����L}l~����[��ć��Ȩ��c�ܿ6y���d��Jpf��tʂ�2c�WԬq�Jp0�_J�`�i��)HI?�A��K�#3�G�V��q�J�1�#��#ƽ>8	2a�J#�l,O��Ү�i��3Es���=»��6�2Qe�3���`ޣ�Q�_�,��~\8�RtD���m˳s:��D�.��K�T����6��Nh@���5;��i����Ur>�໔�;Q)%��~Pʞ�`�bS�S��[�C�SU�fYީ:��_�7����c�iI�2��J�r ���:���,M�!Zp L�c��T����dء�|��d���D�mY�o¸��ba �y�D�		[GP�7�x5YI'X�6������#����Py N���h���lZ]�H�-���3��7�O$~����I�r-�[ ��&YD�	O��w%�����Df����8�'�D4^��C���n���{ :4m}���7���_�]
uN�פ�P�]�c��������0�KmІF���u�C��6M਽KRw���ځbp�ta��[�����+=r�m���F��|�x�ug���$r�y��Q'���w�ަ�g&�O���$�l	�̒w��y��7P�D-je�hh�c|�\���GE�.
���*;V�l9���.�_R�����.�sD�.W�L%�'�9�̹'��U����7Fd�갪�j����Ё<��m,Yl�Ը�g�ع��ˑ~Q��j��`9�ar%;�0��u�iTܢ%���2��|��9P��jgml��W)�+���F��b�T29���X��8:�h��Pk���3Y���ˋ鋜6ZP�kg��8���)��P�GM��z�}�*U�Ĵ|��^���ly ��k}iWd�{��LR�.��(�k2���r���0����G�:}!�#Jwo�3xHԮ�6����`S�m�N�"+�|	a�= ԫ����%}`�wi�cF6s|^jG�l�h���¦���L(z�4DYP���b�Ǆg)�H���|�i�_T����y�����_,�bs�^d9�;��ѮE;S����K�iZ8cq�?CÄ�!��?j�����X8�������{���(z�����U;e�z]�C�fl�� �U�.��<y˹`�͛����w+ӗ�2.�p(}�;�c2�;�,	-�0���r�Fl_Cj���������V���'1��ß�61�S�i2a���=�n'���mgz�&e���m� Ɉ�]:(�f�f�^���ş�Dx1ȩWk�:��Tv���@)���Oq��6o�X.�	���	�gZ>H:|��j��	!<� �^����j���x��<'91�#�|�,���H��=U�r�H�"Ť�d��p{C�⺸SͶ#9;2�E�
�����уpkk��>*:�KĹ��3M~◜�O�m��A�V��0��@%"~n���%ԃ�+P��;_��i�`f�)�����$���s{��a(����v�7iTj�~Y����Ϧ��X�>�?!9�Jf)޵�I�����΅��+�%�1��J 𺲺t�����a|k����m���RMh����؄��ȶ}Rh�K�V�A��+\à4�&Y9���ޑ	�S�X?�D�����G���ѐ&��ں�S/��-o�$�q���A[^�_�s�cmw��O�]q(�������b�+�I2D��*K.�Z�Fp�+�Ǣ�f���
q����$h��B�v�UQ	��_�@�S&؅n ��#�4*�؊��� ����DA([Lc��Ɇ��f��"�����S�!c���Cv{�agn9�H�= ����${C�v�߽�s,\��T���%��\-�j�c2����\4?�1�ML�_��G-�|eSfHo���6|[/��Y�q^��0n2��5�<5쏀�%��O��r���/�Ժ|6���)�>�P���&�Sx<�k}C��C@"�_P�4*@JG�{�*¼$����Е�1�el�(��&��H�US��	�~6D\�w򦀾|�T�0���(-Tf���@J�:����³c��ʴ'�$_ū\O���޷<�O&k�:���cg�oF��dhێ`��L��g4rQ:����Ψ�%CD��Q�q�G���l�h��$~�(�E��]\�IZ��_��NĀք��Q4�M^j���2�=��Z�6����=�gk|�)�J]F�zt=���MU/B1 eBv�#��#�Z��9T��9Ob�N��:�JQY4D���&��D���X�FA���J|P���5�S�S�j��A����&�֭�RW>�D� �D�%`D����O���x�[��R��\r4o�
X��AY�/o#Iٶ.�E�]��D��0���$�Ҫ��tC��6*J'B��*��e�.E+}|�s����t��U67I��4�����ڶ��A$��N'�z�;Fd�{�[����#�';� � A��y�r�pK�uV�(��f�r���V�i�^��L$g�>m�&Hq�����Z����a}�Ʌ��������Nf�O wOʲ�#z��:���$��I�P!�M!��wq��v)�j���E�@�ITylm?S,�����s,��\ �EO���1�v:��Ej*>��&��`��+�AH@A*���<��		�L�q�e���u��u]i��F��Il�t@�� cd��^n�)��5l�
�o���s�Wac��_��N��<#ڇъa��%���Kn��Kd=�{���L�F�Z�ò�J%�ŃM��F2��RGK��+N��s�eA#�s�-F��H�7��Cj�`8#�WGD��q%�S&�������K����;g�!�	�-�z�}�(�3ר���G�-G���_ �|0,#CL��G P���K0n6�=*���b�-<�Ĵ���4�=�Ja�7�Ԥ�/���?u8��B��I��>���p�z�y�v���8UkU�w�H�@�6޳��Nm���Sh� ��,���Ͷ���_g!�Yp��p{��`��b�u�͟��P�KDr�i����
�Y\��g�	q�^�c��1��S�����<K����L��̖=[t�e'�>����r� lh��M�cǮ�����U+b��d&�a��@��c�Z���K��܂�dt5c�2^by��(��
 ֡*��R��6��L"���-�M�˔��Cv�z��ɾλiK%������4�9B��Sqs�Q��b�Q~SKMb_e��*Ƙz7>��Ջ��M����[�c�
e��b�A�����(������z�);w�~+��(�s4G��W��` ���JO��s7� �i��H'����){8肷� 1�	��B�.ӽ�3�������X�r�XQ�?�d��s������_�=_C�1;r�-P�n�Mꡤv��_����b�M3��a�	���p���j}ƿNh-�M�|vH{d�I�����9Q5�����>̤�޿ǔmɖ+r]���R��7L��A�Md��R�c��F��!��(Gb�&6E\��H��������H�Y2E�n���m�_y�l�S��x�	��Q�a�!��(Ј�ns�%S��m��.&rŎ�߶���0���KŖ=�U�� r���G0Y�����1^������N�w���Ua��o���s�:.�~�tL|���٫Fn���K���LV�l�����L�U��"�c�i~\.�I=�<�$��ֳ2���Eo� +�WJX�2�褽��f�H��7������PP��<���B����`�_z���Be��?�8��r�b��q�����Ev��$4�C�S|޺z�E�"�מ�ę��\����E��3]*�
���W�	gҚi�<�yZ.*�,�uOqp��4Ni8_�F�\�9�ۿ��*��*n����+��M�G
���H�3��h��t����
�����"f��!i�	��f#��<zp�aІ�J�분�1|����ʾ`w&����
 .�(	,B.�@�hW��R锲B�� [[x�.q��+%vo�m����P;�X�2�:��fC���W/��xx-@�:sw�hT�Ƥ���i��Z�P!�(���OL��q�tAm��#H��v�ꯚ
?�SV4��w*�Ӈ��wgf���V)�����^���]��ǂ�h
8�3Lm�
��(�DGa�����Y�	����<�"��[|����l�:?�^��zӕ�H�B��2��]�������X�4�<A����ƿ|Mܤb�g3V�uN-1������`���~�LV7�G�|Vc�əHYh5����1P��Y���n���y/�<1SG��<%��dc)
���<e�%�ךS���O=K�i�Gn�dT�w'Y-�g?�}Qb7/��ބm�"6����f	�A/��iZ?[	�����PW���Ɗz�X������>�0O�8��B�+���zM��q9�?�ܚߧӻǖ��q�������� �]F����F�����-j�8�l��	�7k��Tf��G�J+@dS�E��m#��,��[{o�g�@%����x�0'SAI�,�������u�"Wf��V��8��s����!�q	T	�FE��C�a!r��C]��~��
}U��X,
x�{��T
\ha	 ���"��W_��Ucv���-̚�D!�uӲ�����,�{/�8���a�Ƌ��a��qR*���<eAqS�Q���<,�ټ��C�JH�ꔭ��3�&*�y|Y�X�w �nv�� 
'?�����h�މ����U[
���+8o�+F�w5p�6�o��R�� ��M�X��[��⫽�68K ��'���J68qQ���[e\K�pə��j���(���SnӀN��Zȓb`ͺ��+��_�;U�j���������z�2��/�./�袖7v�3w:{�Qi �F��g�,���@�뀱�h2�ꞣa�KP�BT����*e{H�ѧc�c���-�=x��
���C2�M��¤�7�To��V��p��b �]��E�F�+>����ǅ��,���<ҫ<��Yq�
����1��sqc)VlU���a�3��
d���Fdu��6��y�av��,}|���:/Ze,�L�Y2�S��Rѳ43�����-���c��s�ȏd(({$� �6�|G��m��;-5�"\�B;�Ƌ��KG����׻���;b��ޭ���<u�+I���h�PD��M�(T�m��@\_8�qN
EX���㾣�1�1C��G���j�P��0���EX�A�G���!���l8���L�E��6��]�)��e�&ª������q�Y��x�f���Rȶ�e0�1��/��SNh.;Q>�t�+n�+��罁�B�q|Pv2k�j�)�jc�fD���|�Q�#�B���Au}�tJ�7�`>Nd9�4.�hlwL�F�bR�*�j%a(���;�`�� �hX�����6��%:��	
2N:��]�����~5)f��@9���\߾*�%u��q���1��s�(� ���&t�l? �5��5$�cU<��-ǦC'��lp4��W/C�
�I�Ð�sg7�>P}� �!jSA	@z�i�E�3/���AF⺝�)W |�T�߭��d�&PZ�Q N}�\�6���\>y)�lȘ9�0�dЩ�E�0F�z!k���J]U��ǻI����>�@q{?�f��
O`���f,᛻�Ft	JZ�9����,�OpQC�j�(�=����>3V��V�`���%+�pv��8���J��(q/�-d���o$�+Kf��>�3N|R����7^X�EJ��.��5\�9���[� �7���pS���`�ʛ/�P=B��a�����c��0��-�#y"�9�� %ثҗ�) �A6�Gx�=��=��;"/-��U��y�#r> OW�!}�:���]
�����8����=B�
~ǙT$�/��	����;'N�Ū�{d��b��ףz}��Vt˯�Ѻ3��he!���5���_��@܂g�4S���F��$�+�o�ƌq��������:��u����P��h�u�$���w����l�D��oN�P��	Y*��,��﫭o_�s8����Q��A@�+�V�$c�-�!�m���&�/7�vN.�^9xvRj.��Dȉ"_�[W�����@��+W� �/!N"��&,q�^���5��rނ���?�4�{�Oݶu��N2KuUsÈ�bvE��G�+p�9�_S\�i^Ki3��׶�PT��Tz�~�K���0&��X�j��}_?�U�|�X�.��Ū�h�����?���{��7����
%njr�0�r)k�˚��"��6�|��h�Ay�j��Ň`qq*����|���3Ѓ����a�gx�&��$���s���f�B����-z�n�v7rvĤ���
-�"Ɋ�X�,����K�s'��6��`֫�
X���dLJ*;���~6��u�V���g�^�2�������'��S1(��G�=7�	�	�I�Y��^�C2�pхG�2:��Sv{ޫv�'�_�v�w�	������2� � C^�ZG,�m��誁l$.�����t��ω�X�XڏO)�x�%pa}�L��0�hE�A~��"�ǐӿ~�]\a����`��2��ߚ��w�b��}ߑR<�g!D��	�]=ܵ��e�޲�`�	�V��^�����@亽<��X�`�J�3���,��t�����v���7��k�J95�k"��K��y}�"�-c�-h[�WIz�T�]�eu�&ȩ�`K�DU������;�s��x3�x|�x�䞼�<�}dp_5�NwrV���	���S�����{P,/�R_��B��zgt>y��O�nfy�s.��{u�x5�����%bt��"�:y���S�]���_����g�b~۽1�Db�4��!�J��������c��ǐ�S�����2t8<$�G��'k����Q���M��Kv]��_�,G*������/N|Ҥ�ԂHW��+�z��lB�w!�,�F��w|����̴,��!$�T��ҋ��f2F�mqĈbkν����}����&�8�"(��iqN0Ȭ~��H���I���<.���8yD���|����9ѡV��&GX���&��֞�K��.O�A�{��T���C'�>_6�-�_��a��喹{6{"6�����XѸ	��GF�O��w<�:e|@�z�9%ۢ�wG%ٱN㘫�cM\3l��S6W\����@�������� §؂!k�XrF_���s��C�"_�hJ�"��$����8�N��/�NO�Bn�̑�x
v��ͯ	�,M���@6��Y*5 ��Q��tb��9[p�|�_I��]��4�Y/�l�3�{��!ӟ�|UU`[�٪"��|�Y �'@�_��8�`�V
����\��`tdA��b��:kOF����4�z�;��6o(�d<+LRdqb���XX�>zw�uLNy��֟tʥ��1�в��6H��l���zc[堫{]	>�u��S�3F���wO�c��U4iԂ�(��m��{`��?�.a9X�]��rC���^����~�^�Zױ�� ���棁�5���1�G������F)e|��>�3�t��E�SI�6����R1OM���IA�uB��u�3�^�~`B��/�m�'����U��L���\�nU^D��i?j�%�'��W�u�,�Ț��Y�F?�$Bc�,	��∂���7
�hwy`,�p?��>�Æ|cx��OX��
=~�!�v�8�Xj�?�%��VF�e��S[��]���ٱr��f��R+6���(�~�za�x(fcLTa�V:-Ʋpwc�
O����"᧵�P���o�r�/�?���, Y9LU���<F5��ܮL!�*|�1i�g��J��q8�-�B�0�L�Iآ����y��$���/��tbO6�"����u��t{��W��-#F�����o��U��B���͇4�1���;Q2�Ph,���q>,Թ��Wx�.^	f�u+k��c�l�������A�������Ag�af��$5[��ўX��R���{��\�F!�uíw{[/ןE�v:�'����r�_��?&$#~9����i�f��[��b��8�j�iذǬ���S��J���h�Ӣu�� I`�Hv����Sl�C4�g{�2�Y�������E�֗�2�Lfi��U�%ʶ���D^�ięȴ*��G*�l����W�z=a��k�nl�N�}(}������a�o��mpO/���X/ihg�V*6�0����J ��1-�l,��5V��V��8jI�>�d5�4�v9�=�>y�����ʡ��&O%�~�� ��k�6��af(�g�b� H�P���[�ڂ���C� <����:;Q�.�#���������Y�!i;�ףo�ͦ{b�&*�.��e%��ak�W@�P4J�H^7-����	��|p��� @��!����u����9�8�g$��Z�XV/W-�=1j�G����Qc9��j�o��8�o��PD�>�I�G��ۍ�����Ռ_�5|���9��$�EÈ:Z���[��^��/�@�/Iˣ�
�Ά�ac�GW�K�KD"ڰ%�=��T���'�o�5�׮(���P̚�]�kb� W?�#g߭7�M3JL�0Eҿ���x'�K'F����(n���\��I��;c��S�'� g��]��Z�l���Ln%�.x,	b���ߊ.ǚ ZN-�������:4�T��3�c���t�3>,І�Ĥ�Ɛ�J2f�V'�]����y'��^#	�a2y�N�� ���AP�g���f[�w/���3V�+���_*hH�YYz'�c͆�v;�/� #n$U���&���w�q:�.Z4��yҴ+�m�r�a�Bc]E��@>�u�}��^B޺���D���VSd����}#S���_uz#�?�H��,nPz�`O!��T�,ܪWg�8l���6������V��WNi$�ח��%�U�_b/��,5��g�D�
퍰�ttP�h��	l�;����w}�)�?�$��e�$��zZy��-��>�1�	�����aPթ�R�u���P�#�g.���q�h1�α[y�h�榋���0�s$F��2��	>��QE)n�+�j6�HJ6�FT!��X��_C�<ڪ����-5��Ŭ����?�i���GYݨ�kɹ�� ��g.0�n�.@H`���b-%Tߕ�om��MH\ ��6�^�G7�sbd�]���/o��y]$�;]����ls�.�3T�d�焃�o?4XCp��k���� �%��:f��Ц����C�P�"���z����7�\���j<��O�pP2�����
2���s �2��"�R�q��qH'$�op�G���r�N|���a	֩˜�F��^�"bK�i�j%�=�$&[�;	�����f;��y�h#yɾ!��_��*l7f�!E1w9b�G^�w�d�e0�c�\b�Z&�+�$k���/K2՚���2b5@�LK�e�ܻF���0oXJ�e�C��q�{5p��z�L�C��0��+`�p�;�z��D�<�NtB����������
�RT��)L��[�S�,dۖ�H�� � ����#� 7�f7�p�� ����x�>�蓌'�E9g�l�+��g6������~�����އ@v�7�0� ;���oK���ܑE����w	9E)Wn���?S.r<?���>�z2Q@|2yƯq)��=DݙOu�����/-t�L�� yk��M��U��������
V�c��^���s����D)��6[̒K���^�g,�CR����4C�o��7��evk7�؀F�ݼY�99�ғjFgD����͇J j��{�_;��%@�c��S�]���o����$��{/��dc{�1�ޚ3A�BE�����,�S#��qYFv_Z)Lh.2w.G��y����� �)�.*���\��G��
Z��r�МC}>�ȺǙ���s�!7����,���[��t�2Y+�3�ˠ_���b��9>��$T`އ~��<XuM�_d]&~w[��7�[b��h�};S9k��7�����V<��I�j�n��4�~�+W4�`�^�����=G歭S�z�v�[OV��|n���Rh�e�/�o�{��REwu�|m�
g;�c����_�w��r�ق�<z��.�"��XF(=ȭ�bW`���x�tK^����ý�7�����3��ۥ�.�}ptEA2m|���'����S��p�7+�&�u��/�d\6lNJ>(>�[�F9��Xǎ�:�Ҕ��нzR;sGqL�>*�y'T�ݟ�$�����i\�����T�^6+>�9枃rZ&�Ru9�}���޽4��4��筊.�u�LNr��7#���%@D��br���|��tn!�%lAtRȎ�u�4�o��քr9'R�e���u��G���C��</��i��6e�O�5sp4�#z���F�4�U�c������,��*lh�q�T���"trsN����5źg7W�	Kq|ӸHN��P��\H��Q"�Z�x��Z�Ã H��"]wl��;^!^U��c#l�_���z�`�vLr�����eQ3�L�������Ǐ6�0�}ٹ��g�~G�	n%��Gu�X0�-W%�)t����Y���&��18|��u�O��I6Ḟ1��/G�]*'�Ѭ��?,Qk}K��To��W�{.^���;]�:�E.:Y�{k��6�#O�z�A��J���l�1ƒ)pfdǧ6o�����J�۴.�?0v|���ż3pD�&�${k<&�*����3Z�&9��.�'ʸU��`�����ˁJ���e�CN�;P�XCn���qe��8JeW��:�	(CZ�a�͝-��|O}?���sAaQ�R��vH>�8Q^*TrN1��E�%�nA�����=���Lð
渌����[`bꬭuS�����@l�t'��t�tv����oI�F|s='=!���� �=���h���'��I
&ox=��"N!�K�U���u<���3b����=�1��rk���("�aPC�#7[�R7� ��LOy��'ߌ�P�ׁ<�E�;�N�po�,y2��w;Meow����+\i���G�7���RW`��+V���ʣ�Ji+ߦ��c~h�?�e*�4ZI4)���TY����X��}O> �b���>DF�����Z�&�§ݻ�s�D���A����0�r�G���Y�44�D�ܪRT���`C�a���f�5��t,Z��ርYP�\ٿ��
�c�Z��c��|�6�"� �^��L�]���Hយ�$c�^����
���/R2%ޝsټyd1b'��}G�:������P}�(
�O%�8�#mh���4F�ͦ߭��%ru��s}�*�묎G%����f�|�Z}m���������b5!�L~�gZ�	�k甊��o�&�m��<
���@�M [����#���Bm�P��E ���U�����t8�N���G�'.�UҒ���<]ʚ!���4�E�N�r��T�9#���1;�M-��'��&�q����O(��Tq�ƥ;·P) b1_r��gƱm�jP�H��9Hx�� Au�_��$˄^�0��٨�R���	�������;�8�WW�V&.c3�%�7b�15��$�k�oy8���絏��wC����h`*n-|���k�&��::�B�#z;�w�~����F�׎�����dti�����`�A"8��ߦ���w��I��ɚ�-']�bj��X2��۩T�-0������ �����&���^d?�;6��*���f���G�M~V��^��F2#T�ю��b�����}4������Z�loOO�Q�7xf�7��3��Bf�uk�n𚶋cŹ�����PH�(gG��b��.s����I�&�ajh�D`�g����I�P��1[W��r�7*��\���aՇ��C��j�ƫ��k݉��U%"�K��y���㬙��#�x�c���.�>gL�<�ķ�?��^���-6���<�7Q��Z�uz$7̢&�̳�CF���M���ӛ���Dµ��uy���(�Q���a���ӰXkG��h��r�����C{x7�Z�����2��ɚLh%)G1����Nq�+��Wm������]�!�I��M�z��tC*�����X����J�������]D*�qBO*7Ĵ�X�>Q�֚�m�*,ko0�n���i��=�%���t�m�l�^Je���}�*D99�� ���+��F1o�0E��m
$@ �Z'�we��R�E��7��h��5.�@���r ��	�q���������#ۙ���?W>�&�tV�>��T�S���Y��'�|;Vk*����l����ϝ;|<8aQ$>C�C��7U5�@���d��j>3���i(Y�H�#���@���G��E<��L7�p����,�[��/���ǡ6��U�y��Tt�g˽�|#<>�Hc��z�Ɛ�����lR����z�'�I�!T�F�vm"O������N?�qA�[�$�֊��>pq�u�D4��Zr^�dI4B�\�2��YvܻsUY��~���\Fj���vխ����эJ�5�BqN's�S�NO:�Z >�� R(���+t��'���t�5领G}��4��j�×��h�$^U�Al�s��V�i5��u	�V��;����@B��x��+�{��@�)*vS�qX��1hy���(#8fhh_-"�RdeUI�A�~� ?@�d�k{;q�E:ϊg�*%�'rܲ=�H*Z)�|PuR��Jy��ђ]@�R��`�Fm�/
�b���-c|��+%JQ�RW%hS�,,���1u�:�O�>G�t==D(LKKζ@�R�a'Օc��[��+s*f�����_Q`��2��T�fI�L����l�:Ҵ���N�2�	ͺ�����
}��(h��Qa���H���㕒��bn'��k�W֕ ��C�����Jٲ��:���}�^�qa��ֈғ�ߩ�F��"o\p��l��c�u˂��"���
��W>(�ݱ+�J�q#w9�{-�KA�~�3�/l�H���ΌÃ̕,8��Olᙒ����RZ9�4�IY�S�k�b����j˼����TU��|#4�����N�>z"m.Ի�;4�:q����W�jS1�Ñ�z����5?w�Z��8�Õ�k[v��c�#�����@����">t���o燫�9�ր=�����~?�Q�
�*�BH��5H��|	=1l���vkI�gŀ�����
g;7 �����?GۡZ,�uG ����s��	'oʆ�g���W���4'���ڗ�U�Z3ɮ[ݳDwU����Z��Ě�n����*;��/9�7��~��Q]��4E{�A��:��DCG��%\c�W����,:B����15-��`k����6����gǔ<:�ƴ�V᫭k[��B�������<�V�{�&�|�N����I�E���:!s��0�B�9$Ү����m	�i��%�ǻw菎!�vC��X4���W�D�]�e�3._ECf"?�O*�v;X��r�w/�C3�(Q̂-J�9P\,V� E
�op~���L�,��w��1��]MR��[	�ąաp���B��h�gjc5��٧��7�ڗ9u��z��/p��q�c-�R�)�U$���n��٬����x���j�Iu�V'��� �m	u��dQ��j�Ag������H�\|La!}b/f�T/�0?ݍǪ��Ԃ;(͘��A� %i��_[��L���W�����ד�n��B�
�z	g����b ����.��_�S�4�tN6��9L>T�K�� ��n��^�4"�6�S��@+��b�t�\Z蹂=z���Ƽ�\� z�E�ٱO%H��QgR?Κ��c��K�H0�{%9r���h���Yۈ��R�����v����V�j�i�����W��32�d_��6�O6��YX��j���+y9c$*`�ߡ�ɹp��yc���=a�i��ct�0��&�ME��4O�%M�`�"02z�����-�Yk�NW$X���E�&$5؋�@l��ġ��|��+~<*s�w�`I��;��R�R���KZyN�ԭ��/A;`lJ
�-$N��c���O�صe+��pmWΘ����lxx��)�O!<d�S�� ���h�f��v zB�l��s�h匛�'K!-��������z|R�����	qon��@��]U�w\@k���{��,����ujݤ���3ǜH"�L��X�X��������Mv+]=$�8spo>ж�Z�\��Yp���G�X��g6w%��9BJ$�v�a��-���-�
,���/x:d������%>e�$��ǉ`�$�9�Ўi/ �g��l�7�Aiu80~��ٕ��"��f+�����@�Ϯq��\�3eV̕�n�a����+}�g��J]f7�����e;t�c]��SWcuN-����i�E6C��g�nR�eZ�Zy��'�\.��I%>��Ǚ@��-n}����;J��Y9�]��Y������PK�)����Dd�[�ɣb os�x������ʹJ�w�����A0�j$2#.�+�z�t��@>߄C1P��6�ɫq�q��@��#�i���
�#�=�xb��E�qц6���4�w<d�+�W]��]�/�,�zsg��Ma��Ҥ�m�*������M/����ƲHuc��P������K��.mH���3��UY��M�"]'4F�CW�G,�W6t`�-�ݕ�N���?i֍݄�F'r��������<�F���w��=�(��rh5��,�{V�Q��7u	��A�"0f��AlZ��
t���o%}���J&b%�ga��V��?\������LD5U�
��@k��M�/��bS�1���\�vg)����D�Ҍ�&`�U~��-��\\����b�- 7QYӥw��N� �mF&TJSY?\��L�s�S���Ѝf�p��#��\?����@��i�A	$bch:)���(y�||�j�}w�U��,$��Ǜ4��]��x� �Q��xTJ>��!3��_�;��e������si�2����m�+�t6�}+�ѧ�_�+~.rzQ��Fx� NH��)�e��������p�p0!�׎�E%J���g:e����{�"p	��u�H{��㚊Q�&7���EP��St�\��}-�1�I���)��>mYf��`�-�׶
�yn{h�ם#c&�AL������b��t�{셗���^��Bêr�9�q���?������k$&�3��4���w�'��M9�Uo��ٸg��pJ{���#]��}��iS��Rc�G���f�� �d��hp� ���C<�����<-�����~H��p>�,��>Jo�	4�P<�x�#nX��e5�U�{0y�G�Q}�'�4��ZA(	�c�� �m�ޤ���.�� :S�0]���`ɞ�M����\e-g��I�"�9��#k�yC�"���dX�@f4��ȶk%0����sh�&#x2�$ޚ��I���l��Mۻ�!	���3R�"������%RWq�h8�͝�po܈��X;����^ʤ����:�´��J~��
����� ۖ��̆Ņub~�ǠKZ�<�����'0���h�H��i��h���G�Y��u�Ӱ6�´����8,t��k@E�(�ʶ^ν,D�^2zϼq������~M���'2�+�����E��~���N�� ��j�/���$��_Yr1��77r.�IE]��ə�L(naV7Ʋ�j8r�y6&��q�A��W���������{'.�`6?3�v}:R�[�r議u����)b���3�0���q\V�xu�;�Zv�&�C"�tݥ]��,�y�{��|����DDkM�W{)���9��c�א����ʇ�		�s��3��kg�-���)u:t�0��<ttһ%�|�������_=rY�6F�(=(���5J)�*oO/�����)�A,����S��X�Mu��HJ��~�^G�{�8�얣��
�U��"��
�v��Œ��>�jW+�9-��=o.�(th�K��Eh��h�����E��u
�q���4�
�w)}���?�4����$um�7`t!����=��iP�DYWoHM�;m��i�
m��>H�B�Ϣ�N�x�D�?6]X���{��`*�)�b�c�Y��#ӨSWd�Χ!�mv��Q,�&�����Y��sP����S���Z`s�p]��j@�v� �8����?�b��R�KP"���@]6��D���\�ЦhCL�W���i���
yw�al�۴�s#�x� P�DP	@�	��"�
�ł����U��F�Z�����%�>����7�P�mσ�ҽ��<�b>���3�2 c�ɩ�����Ɉ���&`�teK�m*=d��Y���?��_3�N���a�'�N���q.�����Ou��6�Fhˌ����hl�[�%TR��=1Q��F}�����Rj�]P�Z�>���Q���쐌�q�u�>4#5D�~����2-GOt�Ċ��CH)�E����T�̄�~�p�&��&\2ư�>��D/������A�#�A @��܊l�q�DH�>%�C	�i��qj�rr1�=�8U�X OP��:�o�Ch�b�7.~)�O��T�z��y��N�y���'�8?i�[vf�&���0�yBc]���l���B�r~S�0��=q��8�o�sɗ ��9�q��{?ku��;����C���+z�}S��() f�qi�
8*�
���N����	5����;x�-\;o�ࡗ}��{Hp�k�N�1Ϗ���	&��
���'�Vc���~�=K����R�<"5Y�5��\¸a���:5Yȝ��y��� ��/��^�|p9	�'~�F��/������i��:=,��Rp���+0�����,�h�\�:�H���8��v!ɖ^�;�lD���oo�{�u������kOFv0[Q�z��2��;��I<!�Ϯ�&U�B8x��>�`x��l�{m��W����H�L��tP��{�!�AO�����B����%
�j�$śII��ʇR��qR�ome�v�H7i�S�R�0S�����Vj�᠐�l��zo7��]=�{�O"!3�y�>?I���I=\.�� ���*rk��3����7���?�ҸU
&U��yu˩$5fT�z8Ɔ�����9��c��y\�	��Fʇ�ˡ������L�������Uq9Ǹ��d�A^�]T�\a�[���H��6/a�?�j�f/��1�w�I��$�̒�jhC�"��%~[�	ۃ�S�Iz�p4M�';ءg0$�6��Qn��I��2d�	���['V���$�F��:���	G��DL��3�5n��$��6^P��aK�������CF~D��Z�_�c����/W����z��θ��K������C�Ta.�Tʕ�$q�slv���+���'@X�R�f�����w���9	�	�W[ν�1�y���󮺻��)[���d\�/�) 	�a^�YX��e��U��>��E��w��4᳉OS{�(||[���ЮdPs�[�y��q\vr:����0�1ɷ&,d��Ѭ���o� ���2�����^J2���"L�ܘu�n��<HY֜7�s|��������4C_#Řڒ�V�d�n���9�C^��̍���qq��"�h�PŒZ�O�����&��ڙy�Ȫw�"u5�h���p�ec��^cm ӆ\�Q��F���ЯL�AO��{�BJ43�p�g�b��-�����r�r�e���!w�<�52�|͹-��ml9 ivE8��i��x�Ba�x�c^vd�P��ѐ����6�O�j��g4�z�\րµh�FŇ��)])�S��~������P��J��<���.�d��a�����*H����߳l��(r�2��7��ZU��H�1x����$��I�s�[ڇ��'�C&,��]}�Ց��"�0�%�D@""���v���4���s=%�;�_�!�j�"ͺ�],ۮ����vb�/r��R�H��-f:m� �}T_?��	!�f��!��x M+������&��hG �br:>ε�j��(�H���g�v��d�����������T��b���a�楕���f��_~z}���b�\|�9����H�&S���ߟ�3'$�%M���𝦗DJ�>eH�`�os�oR���r]�AQW�,W1��0��)�AC���}�.ƙ]�>�z����'�0'K"��:�ZU@<_��
��%�ڮ�l��hVu�@����2�˶x�]J�V۩8i ���$��K�=�J!�$�2��.��K���qp���J���(�[����}zFv��&ZI�+L�/�����`��n�,K��������"%>Mť�8LR�Gɰ[�$<m�w����P�@g<1P�D��\k�59V<5}�����ۏ``Md&����uu��dη�{�9y�W Z/����B�wD�,ݚ���V>��Q�����g"Qm��M���Q����dC��$X�!eqv�G���b�,*x�K����շ#͋�D@��ǋ�E�ڙL�,p9M�Ve&k�2Q�8	�>Ǧ|�^<a9����.�{��u�Y��{�c6�@�5Q�ZbL���@ r="�8+�RO�P�Ht:���z�\V:L�I�y�7�G����� (��33�����R�@ĉ�D����� �6z���H
%G�8K'@u�PT� ��5/�҇܎T#�"�)ޙ lq�Vvv,e:剒��;��a�(Y�Yh��_Ѧ�`d%��-	Z�E�мpA��E��QRޭ�T�E����x-�x �L+�_/]��Q���K���ŵm/��ӀVtX��$Pb�$��{:. �����C�M-Eu\��n�5"K���z0�1�[ﱻ�R#��-�h���Tu�%za�5�A5g�+㺀�9l�B$�T!��]�*�d�ĸ��&МXP�UJ�ԏ�0�M��:�V^����I�D S�\���9��2�Ui�g�����M�ߡ�esn�͢Ї� �\�+(��rr�A�9����p�p���5�L�UD�RtQ���{��s�傰��5�������	��ఱܞn�f�bquu:��5˞��zZV9��o<��2�)$�3y�1�B�Y��qq�uPeh�xy)j�|8�B�M˖9�#�TV���l�Л��ْK��-�5���8T�Tٮ�-g���?�ػ�DS~��,?b'?t�����3ŵ��J.'�l�U����C��~&M��W��SC����Lm�f|Y@�������Y(��剶�-+hxZ��!�c��Eqc��Z���+��@�-���T�}�9`�۠%�7�9ZW��zw�.�R�5�~[J�V�����m���6���HvG��x��mU�|��քQ�_�jZ�k�߱Wzv8Ln[�r
/M� D����V�_(
����q}aD_���ޢcD<K�l�r��R�c��6��}a����q�&���G�;z��6����fQM$�x����H�)c��*��Hk��m�fV0b���zg�B�WW�L�5-7'��>lSٗ,pi��U�N7����$�d��G��cNCm!�;�~��ȕ�Vk.L�ze?�љ��$�1��B^��h&��%x��b"dHG�4�5�i�c>��1��B�e���9��ew��E�mE���z4Q��Θ,i(�]��s���%���������n���ȕ.U�	��HW�H�$±��2-x�j�J��=��V��o�L6��<~�HO|S�m��Z{�̶�9H�\�d���9(���Ѝm�}N����L�-\��%��^�]�2��?�p2(��*�T��[g[Z����]�'�k.B�ٟ�H:������1���D��N��I�vz���At�XH���չ��W�H�֨�]�2���}p�
f\.8�-}m+��;�e�fE�F�>�]��G�� \����֕i������Y��
�!�D�=v���Nm%~�l��
�H�yеͤ��\3V6��1��Pl�-7�C�?\������3�$>�8���ө�P�k۲������^G� ^�P��N�.[�h��7(�T�?qXy0��J�i+�J��->&�m��A&�&5�O�a�C�A�(jI%Ԛ���}������Xa������o�'�:m?&��%G�g��1 +���
Q�I�R�S�ժ�I��l�fZBH�߱D�q2L!�
̓`��I2:�"��i�/q���9��d���Ȭ�X�O����#��0x)�����-�D���[�=G�t��<Y�pЪu�O?6,B�E{R6���R��ͻ�|�צ�L��%���~נ����C}�F�d����[2z��9߭�~���R��iX��:|!J�V�Ew�m��y�����K������)�Q$4��/�yl8�7����DYu<Z�#�����`��N���O8}z��S�F���D�-Tf0�Tp��, �e.M���XZl��M�}����`�q�lZi����C�4�ktS���s~ϰ��1��,�^�r-�Y���K@�������<���M��i��Gp|�%�I����0w֒���G�<��ɶ�ݳtN�
���@�d�%�S�F�}z����Ŕ=D����q�W��A�mȭ����L�%n��m��eh�u��[ �TO�lW��5�b��C}�k`�u�RB���j��lX@n W֖��t����9�x�,��˂�ɡ��{�vU?|��0W���`4R����R ����6�<6 ���0���*�X�9.���t�d�⵿�D ^�i�*Y��r�ʝ���w��!L;�Ͱ/�n�	J�35a!C����6�~����¿E�}�嵝�ڐģR�zx��t����5��!{�����7�7��{�8�"�[�>%k%�L�n2����� ����h�����U�T*If��s֯oD�NVs�bf&����ԫ�)����0a�Ms�JҊShǩZ%�vk���4������0iɡ^E*Ď�2I!Dط�
��ģe��\�wY	��%�uS��P����t���� ��o,�`eâ��v�Tt�mr6���vMA��;��qX�H�|Ka)d��|Y96Y��֬�.W���S�Ȯ�/ʹ�_��{��U���@)�!�5�5�@�>�`��apEi��>&	������\F�t]Bj�
\eU�.d{����/�U10Ot� �ih�t����j��\'S"bv��_q*r����I�e�Y�Gh�K��w�e����Ⅹ���?�Bj�Eǰj�����~v�����^#|����5�φ-x�g�<&I��Q-���1]�=%�]z��Z�Ηg�Y�|3����7�̵R�:�0�v�a�[1 !L��=��8��>��|�.Ջ%W�s*�^Fpg���7���e�Z��Fح=-����t:YQ����֮�RP�fhP��"�����s �MzYU���f��RS���u���V5�k��_^��U�DقO�_��>�}���cC6�4t��`��^���?�C��!C�����P�ܵSh(��A����b�o�����AoZ��L�M]'���G�9�Jf�Y�.��Ac��O_���Vf`U�W���7|�-��5����x�_U�z���0�N҃�lT#K��cz�~��o+�(;tﾩ}�L���Gn�\|�8X����v�%Hqyդ�@���`D�ȭ�X�.{qW-��:ځl�YR��o�^_dT&���)p�E3�l5��׭Yb��[q�I��@xuE���z܁�Pt�����|����K��vT� E����w���x{zЭ�Ɏ��x���B��f��YT֒^P)U!y�0��3.26����~����K�
���z4Ĺ?����~$�dCiF8cl',<=`ká��~��J����N�hm}�c�[_�I�V+y4�&j�K�`4���e�Y�u�%��QG�E��+aAOUL�^/uz#V?U�7)�C��"�h�l�F�3I=d5�|2RF	oW܅,�\]��c_0�+�π�t�����q���.V�\�x5R��p���<k��!��=Zn�	-���W�aa����l-�p����&%�X�}���ж��fE�{�q�! �db��������E�"Ӹ��1P�A8��j��t���<�	5�o�K�/Jj�)��'�S���`�:p�)4罝@�5�r��e��B��R����|v7�fa�}�3��JR��<�bȦ��e�G�e*p�YeN}�O��"H*��%�ɞ�1�H7j���1�$6m���FBn*�&���|ܖ�����⃈�ͨ��M兇P7�>�cWe!ܕ��]�@��^*�
MXGJb�߽�'��X�oN2�e��x}��27����aŷ{l}�]�IO�#N�筴���|�l��CVyxr��� � V��-���-i9j��Af��>����=��emHX�dk�C��t�*W�M:#5�D�ZB^��)��t>��<����IwP�ݴ�4��$*��/?���R8G������[�4�-��\��&�����9bm�!dL�<�#m�����ސc^�;|'�M��Ĩ�.��[D���죊��d.�,��-����n�MJ�-��r(N�o|����J�]gf&*\>u?�6�:����yt놖w�F#��\�t���c���`��b�h��;J�t��D\vwb�Q��2 y�f�z|���P���S����9�s���A��ô��C����A5��A֯kr8
-� E�=D�hQS��Zq�� �|k-Ҟ�;L���3V�XWy�5:��=�ڴ�C���$�Ңh��avӨ�@�g}CՃ�kafV���j �~M�哛� äH�ȇ-RO��r�04�M9�� &#%��N7�����GlR�P��0�T�o����UR�S���� B�K�� ����D^�����$F�#���11_�-�I?a,��̲����9�B�P��_�o���W�+�Y�DE�<�����u{�`rkJ�T��sDaSʌ"�h��KS�h������E�� �r<�u��qK�o���"o��ȅ)JEl)�(��c��g�5Q����'�YT�$Q[l;U��Ґ�̭W��Z�/��Z~W7�y4�Ն�)f L�K{�"�Hݴ=���'�E�,�ݹ�E�E�Ӧ�@����|�Uٔ�����쪿��~���)�U@ħx�ŕ�i��{lk���Q+����m:�q�2�Z�̆�Y.i�Z���/d�ș�y��{�#=�lh�F�[�q�Q��ZJQ�}�c(�S��]S:�K��n��}�7�A( 5�A�L��(�?���lnH<5 �ͣP"��6��A�(����p|YY�s����,^,�{] Ui�ˆw��/�U#3��$Л1�u�]��6ǐlG���S����]7��C���p���E������� ��]�O
k}���v6�>O��2*��iŭ@d��eB���t^K�v��ҏ)ڬbu��=�lA~��d1c?�ec�g뜔�6�K�m�;��K׸u����`c�� ����mJ`��/mة�����lW\{��6�i~'�*b;��UH�6��d�$*c$��]�y��}ж�C���s���H���(��6j�l�o�0�eŏ�}���z�V>Ţzp���}�3;���Y[���d��΄L��P��Fc>jC�+����+�[�˃��8&[l���qy������V���Iⷎe���n[ۉ[r�}y��p-Ex:�b^!��aK��3j�N�d�s"o��S0��M���=�l�T�u�3G����:ps�tUE��8��_q�H��ObQg����5z�T�*�Z2��1�+irLӁH|ɾ%��I�=�͜-:�۶�['�$�3�9��W�V����"+Xw~��!�`n'!���5�qa�wH���k����d�.�.G���e�w���|:pYf����P���jut}q5�vA�ܼ��$]� ��	�ؗ�vS�"PϑD���GY�DK`�,��ׄ�%�U}�g���Hq7e1������vY�Zs���(j�N�ԫ���ž��!y�����Y��:2k��ot�.�Q�F�P�%�d,W�L}r��b��:���_̰/յS��+tO�u���ُ$A7�.n�X�ig��T�D�"؝]���5�j�K��Ш+���'����1�F�q�sx�����	.�	WV�_�bo"{�Y�ġ<�\,]G-��9�%����-"K!߈��u\�g��m�y��d>�3T�ï �̝/��%�١�CJXŧy�����/��ɾ��
L�M>Gk��o��y͙���{v/�#��d�%�b9�ǅ7.�- r&��Xn���p�e�1�������Am����^	��Ͳ�zk?�;�f:�H�fV��g�tY�,��-�AK�̑�}���G�9*�L~��V�����I�j`�d$<�4�6��-��I�^��~�B�f�f����F>@�%S��ڃ�eDey��Cp{4�~�n�Ԓ�����n0��G�V0�g#|e |�a�k'\KAqL�ѐ➶�,�ya�5���,�/?�+����m6A��i��J�@J�d� ^Q�V���;��|�?l2H��'�qr(��U��2�kW4
Ḡ��!t�K<���ѷY*?��ƕ���,K��M�8��n���s/���yc�:��>TR�=�U��z����-�N����'p���LuĹ���k{)�>�$�o.��^}���������%[�h��2v0c>���Ԭ�֚�)����0_���a�=n�KE�����t�#��9%�ۀ���!u��ϟ�qς>%WrQ$fX�~�h��ts��<~H�??|z��\��k8өjɐ�|�8TXgK��3�5��Ї���ʢ�yΥ���Ңν�c3
�@-NH!Z���8��X�*W�Ns2���#f���$o�cQM���I��w�ٮYAj\��n�FP~�X:;�� >݆��:D�^�?�2����+QdY�Ԧ�-7IPu=0b�bN����s^�C-%���=�]2J�����Qz��+$����b���(D�.��*��J.�Z����i�-ܖt�x{.�~�eg�,��'�� 5�̼gp"���>����
��+�v�b6�or��Y��j�|����D����f���]eix �cd_�(*�3kI5��q���q�����u���a��F����;��q�}���J��-��)(�"2�Mw�<���F�8�Gv(������d�A(3��X�%;q�N�������*X���_]�g��>Ƃ����P#�5�>Ę�)�]0+�E���Gt)�,9��Ԗ7�����C[O����k��9�N����D#�������9Z���꠬���;U=�MǦDh_ֽ��*���\e���Xl�=���c���]��/�_�Hx>��z�������p�,��B�ex��N�"���6��hE����&£��#��[qg��./��`�NTIBе��;�n��8kO5	nk��(>`I?����U/��Z��ĨQ�2$�ψ��V��Y��t�h�\� ���l�*��;:N�#�7)'��f���|A�v�ċ�_z����mh�Ϫb\L�bJ58YyP�����2H�g�f�H��Ò*��Ռ""�^�?�b'��r�R%z{�7zLG�)���*����A��U!���9��
b'9�Y-�Cۚ���\U*+'�Q��z7�]���Y����v�g���4I�%�;IW���`O�y�z"�/n^_�=�;�w����ꘓn�����
��d���8��C�O�.����!^�غ��ɟ_'˨P��K@�����9���[�Lg��m�Q���u#�E �:]q�`Y��a&����ۤ�Yq��Y�?�R*#j9���#4�I��1�b��m�>���; �2J�,p�7���*�[)�2\��Zה ���Ge̎y95x8��3Jse�g��J��_��g�9�X��*��CŠ�2�T ��p�\S$�S��V~�9X�c���_�[.�So��j�]���r�M{����Gm��6P_kŞ���R>sC�+t��nʙ$��c��F
��$  �N�{���)��Y�ǺHC���9u�r
��6V��#�����LY6�=wETnñ�y9��bt&Q����[W��4j�L��8[m��#/�JE>]$P@cjŻ,�L�{��񵵺�e���$Xf��1�@0��+`������	�;V�Ȟ���=F��Wo�(,�#|��+�e���M�?t����n��*V�*�
U�v1���s�`�ƚ���'B�D,��:2O���N��0�E20�vq��_��8��
:z,Q�Q�۟s�c[$:����V�P�
!I��x��4+����m�k�>�tXR��eU��{;Q�zg�O���C���;t�4���W�@��?NPx��:�!,���iw���?ŷ���Y���A�K��������Φ��%�v6Us��M�V��W�	�u��e����z�"<���Z�R
d܇�0�X�)7^a�]��ס���T5KI�(�_;Nȯ�fg�5Uv�����f�)��=ua�|T�ڷhD�!_7%��A<Be������O��-�_q	̂��AlmG�\g$3.l�vw��Ŭ]5M@#��o�+���]����������GH��9�@X\���A�X-*D�����z�knZ�?��UY�k�f�9L`��ț>�`�˸�F�U�{��gw��ŵ�=AZm����X�8O�k��$%r���t%T�9v��o���#����l�9�p���:�I�I��]բ׫�`?a��9Om�ߟmF��.��O�����)��I�2�'9u͆�T�N�x�N,�-x��8��Vɀ�]Kv���!�":�jF���*dҎ��!wê�y۞��c��"��5�"�L��h�Mb�,Y���-[��MĹ�3PL*U�
̟n#Q���5Np0��b���K^���&';4�^a�I��C���f����e�uj�%r��*Ҥ�Ðs��rp�K%̧Q�&y|��}�ZL~Q.���3�,4�0��u�{&��Z���g73��!.�q��A]-�OL݄0����_��3���G�o:�akW-���7.'	��6���MW(�}SU�)������?�z�M^�P��a@z�kM�{�E�<��
���%a�҉�/���ߐ�[0����ۈK
�T�g-EF��{�ۭ���,_E�H�ݹ>�����)R��Y�qK��s��E�5k�>$�������HHF�\�O�Hlq��!4��O�����1�Tۋ\�o �_}g��ʥ$?iP}��@��]L���14�"�%\�FZ�t7-�B�����w��Zӏ�%ά�fi+�����r���h����y2��_j߇'@ɡd�Cc�K�"�OQ�H�[]�r)3�3��	�y�c�PV�B���A�=ayQZ<�����_���2"�LsT��W���k`���"I_<O�c�-̑^@m�,v'��j#� �?ss9��I
��lb3���ѽT�	�S�O�����P��5������ݏX�	33g[]e;��t����eq��{*d�9���iM'Lo��
�
�F6�7G�p�>���B�@��w��h��]��b3~ڼr=/�R����|�4e�x�?l�
�K'��c�N��y(jL
T(�0̽)i���2k�� ��ũ��������_a��m,Gu@���)�`�6F�ym�5ڣ��X\_t~ ��(vn�4d<��5�6ymT�y"���y�zK��WMW�����2@�����Z}j�>�+;+���_��ʩ��!�Yng�U��N1�B�L���.b\���&����IU�Y��j�c�O��f̰�h(<֖����צ������ƽ�Г���f}%@7U
s�`��B�{�dk-x��!��6��:�����@@��;�!�H�h�Szc��YM���A���I�$������\��Z(�N=y���s���$;g��LT���l�*Q��u��^�  �A����Ls�t%�y���}Y�N)Y��� �-�oPY\t�lѣC���L�,�ۦ�_�t����Ȫ^`����t�eBOs�O�$?�v@�9+�5S�[��w�&Dkrf��yK��B��
˧�v���v��"�?���G���Ζ[>FC�z�=���E����(��-��8����4>��6��9Q��Ձ�7ħp��{k�p�T�0R�9l?�Rk�3�4f-H$���[��i�doA�+qw#��M�e�D�9~§SÀ#X}�^;��I����'��u��q�.�T�F�u��KJ�?�eĄ���xʖ\ubԠx�;�C7�!�t�Ǘ(�*��+box��:Jq_ <�ѶG�<�LH��lF�+�%eDիh��o��t���M���ȏЭ�4/�H��+#�L�J�(��,��K�0N:6�8����*ۺ�J���K�1<
~~rSgA=�;3���!�]Z������!F�����C�I^��oes�%�ț�~.vۨ��p����!?f(���ϲ"�����a�����iΨ���o�&��Њ9J�Nw���@WWx��To��N-�l� �Sq��v����[R%����/�R�<���J��*{c4*F��Il!�@8��#Hm���a<E�F���T�K����'��N��ʼSX��V�Jgfe�M5`�b��S�`�٨	�8DM�v��'W�z!	�Ȍ��&�r��uՠ���lS��)BC�دX��f>>�_��WN�]0J���0��vm��W�K�{��{bc��sVL��7����T��X��w6�����0-0i�/x�6�F�gmjL\�u���W�W��s8B���NS|'��ڂ-�R��uq�J[f�N^�o46����ȃ�3]%W�yAKy�*6U�/��I�����;���`6�	�GK���"϶�n���R.�%0�d��~{B�ٓ�7Z �F�ȁr�v��;���qp��_����7�D��(RK�v8�z�pq���Wk,��8H/�Y ���粘�����W��o�Ȑ��y��9ljNb���Z��w@n�9NWm~���l1��&�*�>�&�^jz{dp��0,���\��\�vC�.��^���&�`?�[�J�3u� �x;���������ɝ��˱�A5�L�LA�[jqU=���sY������v�R^�D��/b5wnd�&o�`���,�K7j��e�� o�۳-�	�l��1>d�5}�$۵}�'CX�Z�aQ��!��	��B/����x�w�PT�p-��p�[�oZ�����k��v���D2�����]<L)d~Rh�؆;[��8@�>Zf@q4v�c��O��L"	{��e�FT�:�J? ��N����a»�oɉ�*���P&Q��������8	b"����	����%�=։|�/r�iJ^�2����`��I-��5�pr���>�kT�:�zv^=���$��J}O �QKhbK �pj�h^F9UP�q�*� Ь�ϕœ]_��J\#�b,K�,bB�~-w�U��m�Bfl��>]#� ���7��Sd\2Z�&wPR� ���*Ȏ���<��=��#sȓ/�明q���	����'���`��c�%G�S��X�6�?z���m��L�0�a�h�Q�.w�i��w]�w��!�Ql�[:x��U�E9"�mj��b�ζjge����J��vA����8�*i9/�&ƭ���P0~�%��]eˮFABG�����9��Xn��I�\:�+�jc��K�]=YR�e���TI�t,��(1�1D�U�O[_�������7��]qc��բȧ0��������H�`le��=����M���;������A��������1��-t��c�`��߈���O|�uo� ��;�  �5<+���[%�["�A}�n������G�zF�ܾ0Χ��x2�d�^???����!�3�o�hHbd$�^�e;�]0V���=�0��E:=ӌ!��Et�i(db/B�m�[ѵ�o����U<X��ܣ�p�v%��$[/~c0~y\��,:.���M�o����`��5F,�:p���g�|!�/۫��WۖY�xl�P���N��
��WV�v�	��_���J��L�1G~�$�Z�6H�x_�-�����I;�4�ʡh�(}����� 1n
c��غ��AM��+X�r����s��f�C�x_��w����y�6�l�ů�"#@S�9卞��q8�7��̴�o� fm})0�-k�|��Ղ^�����u�W7��	��.Pҁ����!�N�o��g̟^��~��?=6����d@�=���-�Yd�����+�j����{�"��[�(�B������+�k���N�X�<���o��4"�����^B<�k��O�D|����H���-qs�s�Ԝ#>d�?�Os%m�������0k����y�7��N����[��W�ˑ+�_<f�����p������#�?u�Z�Sv���Y��:�����,�x����f_�a�d%�Ŷ1O	�,��O�I�Q�X�/��5� W,��� 	{�k�Ƈ�	��ٍ
br�1uO=�VG�*�/g�d�	����aٍ����QIֆqѿV�z�ڜ����kut�[�,��)x�ͦy��6���+03("�k�/���z� �X��`&4����%"G�x�M��1�{h��|�.��*J�c+5ϝp6׍92�dLJ�G2��]���+�A�%O�����hi���<�b�-��NM���G�����8P,˿f=L����w�����,������W�Wb�HRB��%�g'��JuG-t*��9���ɃB.Yp�a�W}�^ڠ���,F���e������o�����>��(#�u�}1�6��zfL�-�]�߰>锤)���(I��a8�ٸ�Uxx��]/��=t�-?9�������8e�q[��ݏ�� 4����|��)�>�¿B����# :��)�xp�l�N(����E�e�Dh�ŭ��43�j,�|�*mi�h��T�Nx]>�@p;�k3T��9�Uɨ���Ʊ+GĂ����8�u�kì�l�U�/��׎����;P��Љ���&��X�}f�Wa
86$^�!a�0
����x?��QPVM>|yK�{=�P���^U0��/�a��(��7V<C�a_Š�.��E��zĎ��`�����������)Ӂ%4�G}x�U���h���A�Ks���>�圚W�2#�*�wU�	h�Q�G�����Yg�K��c.��C@��f��1����"5.�]5�n��L�_�5#x�9M�m���ث��'Cm2{�'7Ɯ�j��eb��lO<A\p6��N����(�B@)[���������OJgd �6A,Z��zo�w^����Ww��v���l)4��X螂��]��P	�'w���n����;�����hj���r���J?XxW���ټʾ���i<~��1�g:��\�iq�ݠHbBU��*�mk�.®,v�G��B�ݬ�
K}nRPy�a=�n�\l�z�g�y�v�L$u؟$�{�L��H2S{�E��_�o�%��rW�FR��D�b��£[���p�E����l�Ɇ�*�XĽ?>�J�>�_�����㿳�Bc���\b�ؾk=��Ĉ�"��t�g"q���Aad��9bpc<�|ó��]i:u���(�`( 	ZO���10��B&�~8X��u�����	�`֐z��yMJAFEo�Aly��5"cG� �ӫ+�W��!¾9F�]��H6^��8]w�|�9v0�=�N����X�n��Υw.\�&�\�`���̒*���#�P��No�q&��ҭޘY#0�%��E �dosMD1z ��y�o�&�[���\Q6I*��'��18u�D���6_�|��u�툸�0S5��(%��7Ń�ҧ�mEI�]bQ~��ݏ@�m�6�0`��L���J�(�������R(��.���_�4��&C�o7�e=l+��@צ �HU"\�|Or��@
�+[Y�$$��GA^�@]�8���]I&�3�I���ʑ���E�\=���l3�%����kIq/$��SN�C*_���|��]���yd�� �����M7q�l+�����!�˲�8fp]�$�Q=��a����-C�u���l�V����kRs�V4﹋wU
f�yv�q�'{���sT�8g?�b�w��1�5)�O���š	�,꒑�l(!.��_���d�S�F��zY^���kSx�طo){+��;��	��wJ�x��5�#���&�V�;�6�)������3���BOg\�y
ºp��w�26[Ҫ��E){IÊ!�Ov��6��}xnմR$��0��[X�#�E?��U��HB�j ���W��G�J��>57�.:��bHB<���&C+S5]�R�ۈ����4����Ӻ
�~_}�E��0���]�b��u����$p�]-�9�C��Bl?�5ڲr2+�Ґ�(�! 2έw"W�p�2�9*�By@X9֡x�5�]Pd�N$p´޳��L�����,�g��i�[t��۷�u����`���=��g�DP�]tiI��B�օ�"5�����no5E\yvIҌs!�kk\��ڔ����Mt��h�l��Km�^8�+��q<��_�.�x�Zr� u].p��5��M7�a)�5�D��ȶ�_K+���7��Qh�9F+jɁ�l��'[`������%<)�v�#��b�ֻ}ڐB�*;�V��� mW5뜩r�y\�r��l%��9��n�4�H��i����\�.S�%���i&E
��Jf����Sp��2T�x/���q���?�[,�fp�#:�9.�_萘������&�|4�Qʰt����v�D�_X�L�
��	��*��W���5��Ň���[c���,B��)�5����F)S�L1��k�`�2�Gy{��D�@�d��R�kk���{�ݱ@o����Ӿ4����r�#X�ߛe}�앋Qt����)�vBD�S������z�qŎLRh�J��'7��EdA��6oV�%�ZP�;�<���l�'c?�Ǧͨ�#]�`+@ku�}�is"�RVy�u���M��_��P@	7A4���_]�d�^̪�i�Cf��N�<�v�M�5���.1)���r�7s�mU��(F&�Y`�e]�\�J��c{-�u�HL	�~`�w�'�L���v>���Mޟ�rq<
<Na����zd�IU���b�j�@D=�� ������$u�t������W��d�Ds"b�U�0�\��~���횊�o�+BK0�1����e��>�O#W�t�M�	�����Ĥ�
�-LK�9����	�HJ#���.s�|���	� ��)��4dZ�ϗ7�8F�|K����e���)���>�|��L�6.�%��,�Nu�$���\�K�j�cN~���JRױ[��l� v����Z���Ca�)�2��M\��õv���4��T�WO%���0��(���Q�ۨ�����o���}:�K	�7�L��`���+�lF�K�p jorh`�>�� KB��G1qw�j��(�L ľ��u�:��m�����(Et)e�A)�Hk�%ͣZ���Y��)[%������ ��D��\�o�ű��y�=���.���N:�ه�쮹Fހ� g"钟#9�����c�n��օܺ$_��{x-O�*^3�.?V����� ˗��񣭊��1��F�$
�pE��`��G/��*��	���1�����w5�;v�f���u2%�?Ɋ���V���
�LQD�$�]꾢_y�p�q3���U��ߌ�e#�����䦛T+nWs+ozDR�dܱ��-����6gMחO�����aq�lW�}?��3ռ]f�cն|���Z���U=F ݱ����"� l�P�yf%�/�>������J�����!W�F�/��)��IK�BX>�Z�8٧Yݥb�t70TnD���4�*}����نr�C'b��/���
���Ο//x��'�H�6�U^f�(��9c�o��A�H��H~YקElI>���(K��#��f���]�{D�(B+xf8�����r��3��z��5��H~����Γ�&,=��H�24H��sݢh5�M."�����?�<�=B� �,����P�nvK6V�.���r\zR%X�X��� gG���u�<U�S���5'�Y�D�!8���,e�~��w���T+(��7$3�i�������SZ�� ��#����sBY]��l����^;VV:����{K��Q�i�F���#Χ��"A��{��k�5��O)���W�k���6��\���z2�~��(]���Ь�nh{�i�x�lui4��k����8�;�[���XO��4S�O]��G�Sr�6��2��ʾ��)1�s���LS�n��Q�]P+�PQ��o���R�^q���%^�N_[��Y����\쐍���'��/[�8418ۅ����KI#�/��3,a�}�9P(O���%�9��u�e�Q-�n��� +��x�z�L����rsOC�q%J���!�׀]���f��������þ�K�������I`F�!�q9{��< �Ѻ���Z��7��P�c�zÚ�!F��%K/�����ЊLU/����������f��!�kU�%K����f\?��&�����f���$�ڈ�W2�m����UA/[�<����T���)aW����q�.;��k��rKb;,#`,�Y�Q�S��b�ԴӒr��V�H�Fp��|Հ�8�+W�f��H|�PQ$�-
�M2�Z��]��י��ʝ���$��S�lnYf�>	m�T+ͮ]��,�o���'�h��E)^K�����{�:���A�R��:Nr�\~p�U"g��Ӫ��r�/*���C\��N��Ce�����!�p1kpr�r�v�� n<���@��=��T�/�wwuŵ�$!�F؆����~�r8M������Ie������7æ��7����q�΀�*�?��0�]�$aN�>xG4hU�NgVr�������'�У�I�a�CH�X��Z����N�ʟH`FR.-�b��y��b>�������jDגb�4&�����Z�V�>�=��1�
1B��G����p=�Λ����b���e�OF�kj���i��gt�]�p�Y���0@o���1X.��B�x�ZY��K�x�������4�-�=���$�����/�k�j��ݓ��E�hۂPw��I:���>|�#p_���U� =�A6A j��ߟ����2�����`o]g3�����/i� e2�/�C�� �-L#�tP����%X��ȸ	^ƹ�:}=
I�G�����Ϝم�v������"1Z�B��T
��{V)�0�j�����t�X�{Q�,�ڋls��l7hI��A�2Y�m�e���9�8�%`!�y��Mt5-=܀;���Қ�_�_Ch���R h@q3�@>Nr*3N�r�/�J�W&��Ő��10��[I���H��_�D�`� ������5���p�L�RD�O�9�;��vHt���[p!�'JEH�I;�/���`.7�f�;CԳ�7�+�ѓ�qiM3�-a�E���lc��G�W��{������!�H��O<[�X��_�V��}3e>��gӣr��r]�������x�N���)u�E)����&5U�3�&�Jp]ih�����˥�f"�3��}�K��*�vSxxH��t6�@��$Ӿ��K��8t R��SE�й0���{�V�ꅮ��̊QMb��~=PL�Mlp��Lx�?G����)cbk�t������0���tÅ�Th%� �,�1�;�oUl���F�x$�/�#0����W�DL��9`�C����V�!�)�2�*���(&��&�Kq�5���#�G�)BSȁ�9��mX�ZL}&S��>�d@��l����Z��Vպ����6���}��ʳ�VJ(L$�3=�诪�!���\]%_�R���I@��D��c���u���<��� Y��ֳ�]�Ys�Dh'V�J��áVkPaJ�00��tWY�6��1���l0N{ژ���P;��:�-�V�
6N�o+�sM�-��ųf�"��Z�����C��m���5p��#�^Ik�Ye�P����@UI�~��~x^�s4()N�y�r��2����a'��������z�QŴ��T��es�ЄM����"���C�(dQ�`juZVE���0�!�S_V,��d5<���D���܈	�=����[O#��wa/�qpte>'7ņ�����+�lH��Ӧԍ\zZؑx�-˝���1������6W��Vu��>��]W2ŀH��1ST�����ƨ;���QM#{?Y�u����6�-s�܀a/���qN��X�b�yЃ�&(x2����&�^@Ō}'�&yr+W�-;����O�K�m�d�u=�SJ�H�ѯ��?��s������0MD������D�s�n��<�~�������ic�*�g�hP@���:-����j�����7TaY�4�)����ԯߜ�"�ahnûc���_���č�x�G?r~�M������tC��3����beWOB��U_.M&䶐�P������~�R���3�� ���'<rU�7d;�kI�Ow����{C�0���bU��fFp�:1&�	�^�z�<{���&_��;n�o�����=
�Zi�0/�c�ݣ��ܮ����Q���[�g"�!w��w�O�<)�R3����" ���:�y�娷i��H�N�*ˏ��kF�f�\Mc*QOM\����b"����M�k��8�O3�%r5���������G��K���sM�"��g&�䜱e�j��Lm՗���=��]�`a�Wjױx�z�oŎ�H�Y�� n\*�s�٩��v�O=�/��P?���t�[�'�<HNB"�lj��[y!m�-��[maD�Hr�5�MֆWAn�F,n�j71��9_|,�JpՑI���_N=>�P/�X�:m�~���t^�	<~����+f���������-"��}��������Q�.;P]-&t��<�	?�.o\�>'U�dЎקk<[�@��b7;�Y�1����l�l���� ���^Iy`+#�u�(e�R��t��a|��}΂	�9�Y�K#{о%�`8^��Ni|$��^���c�}3mu�$��!2+.����N�Xߟt(Um0@�z:?�;)K�ߘ�k���LBA0�[�*�Qr/�+���脊�� ��w}���\n�9��Zܽ�F!\^�̺�4�J(�k�'�sQ����h.pY��^���'�`�ͩ�������?���YY\��-�/)�U,�$���ɶ�R9�O$�W6_�#�F��̕�W.��O�~Y]j�,!��2��8h�l�^���×ҏ�>XM@o�X�ٱ�D�l�2���I�����Q�\�k�̭h3�71��F.'G����C�T����1�d	`R��r�ǖ���V������Á�e��.z�,*ci|�
�j�m+Z��K�#�|6Юg�g��.ނ��g�t�js���
�S�U������C�[
����l�7,��?T�L�R�FGy����uJ�H�4�B�͉K��G�B�H>��Z��c$n��*���2"a-�b3��'�M��!�k��!GT��$B�v+��*���%(ș�ȷy���G��&�a�N�����ݦ֨#�s�G�	�@�T�xv]�B��Kh��t��o	�h<F�<��rV5DLr^'� ��J�tGW;X%N�U\t�Dt5RʲQ�G;۾���Ŝ�_��A��-��=��=��QPr�d�w�:im��(ff����g�b��M��J����B�Y�Ȕ/���V$Y/��cNod��	��ʻAζ�O5HI(
&��g�Хj�})V�)��t��$����3l۰��Ы��?W�u�~��k��@r�B���C�]�C��n�K�v4. �c'�����SBcA�?�^B�S��nL����L���/Ѻ5]H<��7�B�'߽-�'S�Ve"��d��k�j������1wN��(�� !Cu���Ag|2��MHY�f�@t����Cr�3�xc��}X�W��H���0��=MչK�7�]t�6�3w.��&�{g�]~��|��N��nJ򅼓��=0��MjO�������F�z�s���%c�3�5a���O���)���[1�{Lk��eߖ����h��	*׵�S���:�Z}x�� �i��:\������d'�fR禭1�`��O��sjm܏�Ʃ�5!UiP<��\��,P1K�5�F.O�l��xnьq�b�GL1��W <��O�k+�=X������l~#p$�7(�
���$է��*Ъ�?��<���hO�2��v��?"Οi<�I�oRv�Zj��!�(���(�"D���۴;�x\��$#�q��Y�����R�@��nL]��l� �ѷ��sk����WB�D��e	���Y/�D�kWza,�^29%����
`���T��6�Z��*bџ��|R���_-~$��ۘw���	l�}��W�Vn����3%J�����D{�@ڙ���#�x�}�>����U��f�n���R���S?��4���=P�.�Ն�9�ΖO������&�Jpbz|�6�*�
�kT|��VH�D����=�#�Pl`�L{��D|G�e��G+����h�g���6��K�-�� >9���w��uX7�YN	�|�^K��lͭ�G�E���L2�����$X�	����l�<�]���}�]��O��>�q_O7�h�a�˄��m@E���m˺te>5%c.�2��V�k���z֞���y�4d�}����a9�}dѰ����s�+�.w��<h���_���n���\{v�\6��3��mE�5Ì5��.OS�$���0�빾�7�,��l^�m3w|�����~]���e����]�uW��~Q��"@"�=$՞`�`�6WB��>Y�@Mb�6���w���R3�DEᣡ=��9�ɉ����=>byAa2v]���'��0�
V:[�fuS��dx��v��ýe7����P�%F�3{x`^ufӾAF�	��r�4�%��k����y�薶'T&�ޡ~ɐ#B���a�t���Cv�5v�[�9�в|t]ә�0��bq���e,1MO�ݺ�� &�U�u}B8F���0�7��5�(H�BkL�@֜�@qaR�WK|OV0�)'�4A}�Vw��X�j�9cnM��E��n�xG�v��49���� ��U�WIl$�MxZ)!X7���>H&G�F�y�i�$�d�Lr��	�d�O�a�W�j!ܾ��BB�8b[��e[�}Be8�{�6���.u��cdHڜO�9yc����|-�hS;�g���in
�s8A�r9(e��9���ӵ�6{�\����W2�K_*���f�w�Qw�9���߆z�9�I���X��� ��!/=D-u��!H/�������):'clāF���������'�S��5��KH.���E��KW�1���.�ga�9��<%�;��h����,�{-�p��;'(A�h�0��\v���Ê���D�}���eN˼�~�8�S��Q��~�54ro�re�s����d�M��7s�t�E\(��P��A]�E���;�`q���/o�Yx�H���}c;A�a�9o4����*��Q�ъ�"�ֽW����:�2�n+x\U�P}1G�)�)�VP$���𭝝75&�ێo6�)�G/�����!�����w^*��{^�:��*Qk+�xu2�W>�h�5�h�@���"zH6$g����������!��y�w��jR����֤�3J��4���ܵ�d�Ci�u��B�����U*�.��o�zy'�:���o�V�7o��C�������l�Ҡ�M1�ߠ��!��ͤ����t.��hQ���Ʌ��t�w��C��sщ������D
Ԕ-`�����U�@��3���c����ܗ�&wn��[�/aA������G��ܐr�qr�B�,�r�^���HT(�-ݓU�_'��͸��T�ǭ�5M��hC� �ޮU�
RDbOg[PhL����v|�J����	Ę����9�my���ga���A,f�����	NC="7���X�	��s��ߋ�:���]�u��-}:�z�=Ex�H�2iY�<���D`$�a�fxNlѠ�7��y�"�?��_�8����>��BƳ52�z�:��)�W��,�d�G#����C'��"E٣���*S~��:�<ek��^ e��� $��8][���~@�F�EX�8~9a�K�^�+6g7�#m:G���'�Po�^��`�?�/X��13*]�Ё�Ky.��,'�|qu��}�=?�U:z3�d�;~��ld3(�ʆ�zf����f4U���Z-t�Q��q�M�偈���A��U��L~ђ�_�a�!]Xۡl��I�%�T���TQ�^��\#\��{%�?E�֐�\����sV�Q�O5yĒ86�BM:1q���w�.J$��NƖ�h_�r^��� eB�~y &uޏwL���2p��V GI��),����F��P�jk�vbK��4��.�"Y���,f{�X� rkIK`�[�������'����nD��s��T�c�;Q���lRF����O��Yv�EK�>��a�!��+$�(X��4EB�4���b�-uH)�eQ
��M�߫�F��/�݈_�È��������'�[��5�u\(�2��E�T��?���L�]�s�Ю��!0x�i����x�9�D����H�q���^A�\�}���M�Z�|��Z�=��r�U4��s.��T��KyoHo[�)����,.����������ir���A�Y%�߃&�}�����iΣ�c��r��V�S}���7f�d�T�
�\ඩήl�V���+�%�Sb��ە��{Aog����z�0=&��x���NTu��-X��i`b���1���^�+J�Yr��yT�H�&�N��[����d�-V�Z�\x�2��N�C�5�r�KT�E�y��a�]�"���P�PF�%��'
�m��O�Y����d���Z@@8��!5�]�$�]ΪaF7�nn&�~S�h ���W�:Y��̉-���Q�^n����FA��}�|�WbP�3�m/�뾠Aw�!��g� m<L�`6����Z�5yմ1���SJ��g��:�i�Ʒ�i�Z��^���~:Ȁ���� Z�L���č��
��Ca�l=\&(���7������ҕ�z��&	��v�YW
��o����̟�(�<皚��KהD�;%�E�,�Ã�����c�����jc�	K�Z��6o{��H���]_V��FEV$2�y-u�
��l�ɟɝc+�s��֤��Kt�ZLh3�d���G���x�w2���H�,�!��"7�I�iL[��6�2�w��' `��yvS�D�O�JI랬!i���5M��F�Ψ��n��9)R��3XD�Ư�&�_ƒ
J�(m ���2j�S�k<N�_�΢"ogű��Z��� �-7�lh������7��X���}�ӛ#ޠ��#��YMB>�Bq(��<'�nG�'tx[�.�c7Hd*'&�6�ϓ}���Xq�7�J=,��~JP��A`^iR섟O��D����}p�}��^�2���#��f��,'�����1y���f�u����vca���hN=Aۑч�Q����q�Os�	�υ��j�aI��j��#\��&e�k�{�q���kN���;�+���i���b�O)�U�DY+H��{��?�'�¥����"����ǳJm �뀲g���|��acXC���>S*��1A%���^0Q��f3�i/�~�Z�i<"ބ�{�AK=��9�ܸk��q�^] �wp*��-%��Ҩ���`c�+2lM���F�ϴ���W�G����x���^۝,[mW��I1@ĽI����h]�{��e��4��i��L0偌��L"����g+���xw����M$t�)1��T��c_(Yٍ����Q��O�$��39�K�Hu��?\F���K�xh^����Bk�T]Ue�HT�2���@��B�y�U+*'�o{�.e�{ڔ[��Lyr����y%�7M��î�F��_D��+��F�Z�Y�ͻE�/_�Α��ƞ^��A��8��	L~%o�uz����(#~�-3�+AD�)^�L�I�O��#�C�/�����c�V����{�o�����e-��(¸����j~�d�5,nԇqf�pM�=@��FO�/����m��8�un���l�Ҏ��%��^�`Q�S�Q)�����Oi%!����J�dD�9��Z� �K���j8t�o�ww�?`�䏸�䊽��=~�3Cc��dT�������}��֧X��j��[5qR�̧��(�ʇXm3XV�ݿ�h��������s'�c� pg����q!~nX�o��ST7�Uc���' =�Xc�/��qm��{�-����L|���n;�%Ӹ����D���U�%�[��j脶S?6�#�`Ҍ����,��AJl8r����e�i��3�ː�6�m'��8?�m�X*Z�߻lJ?��W�z�����8��n7l����k��G5ء�4T"B(�W�rd�_A��1�G�A8�߇K��8Z���F����Z�rn���Ǭ��������I�'�Z���Y�R� %@���,%�P�zws�Ria�A����V(�&��+�+I_8�%�Gz���5���t25�����bWԶ`M�f�t��q��bх�iD�RL���3t\c"&�?�bT�j�iy�;7}(�ț�YSӹ��6f�*� ���HdY��☕ey����]Up�@<�[U�W�%Q�;���n->:'�l4������q�ų4+G�F'�c���5�@���؋|~@#�o\-�-����{�EBx��a�7��4,'@�������r�Kh�жd�lGx:ܭ��A���Z
|ګs���Kgl�nפ�~8��!�Ş��:��LXJ�:7��0��	�>��yv� k�srB6�`�2l}��:�H��#���}�w�U�Z���#��� ���|��#��	�� 6��s�E���\��V�e�կ�yU&A�{{���e��\��R4�h��*,�B
��-��`����]e�_dHl(���N�:c�C)����$��{���T<yfQv=J�� �mt�ց�!�4�0G��SV�(:��m�X_%�[��3DN�*�R,I*d���|��	�6oF�!f�wHE�~&������=�|�wjk�9���o�K2^&�q��;< d�ؼ�Y� T>_Nu���@�b�@�Ŭ��˻L[��B�z���o{��g����
a%�+����O���\g���K��f
G�/��4����(��h���6�$����dg���3�"1p�#|��o;N�ghk$*D'/Z$yUK�f�*1߳�e�_�Μ]��xhX�ަ+@Q8�[�����v�[q��J�&�K}&	�Zs�V����H�FC� /��{�X����:�U���	��yJj/F�Mb�v�.2���������ǭH&>-%�2�������?5*������u�So=�������d���Qp!T�U�m��<����[�^צ��q�w�
���`>������[u��O�s��v��i�ș��)����՟SI}���vx�����ٯ�d���Q��D��f�Y�����h�Lw�v؁���cmK��������1bM6�L���1��Mng ���Ro\�Xh�n�%Mi�Z��׻��T��w��_{6��v=`�S>@5�Z����hJؽ��f�)�����牘~�MB5��'��X&������xTd��hY�N2�櫓 ��ݣ����=��+�!�n�6Mf˯5+]��B���~ �<Ƽu���d�����4�6����_d��9����xY��R�"2?��B,������Y~/�P�Y0�B�4ϸr���%C-G�,>p�f�a�C6��yNL�_p ����M�Ւ2<T�K{����j�s�����hک�",�)���Ҕ��t
)�{Ϧ�����߾��� Q��~EC��YG����S=F(M�f�X��e��.6�rY�b�E����|x!0mJ�;n����^�X�*$�<�_N�ΒK�!(�����'�H��_���?!�0������ �y=]Q>�ֳ�2�3��R��SK�ca��4�*�k�������.���U���f��.9�}Ee�#�|�h��m����}<3?UCkϡ%c��]V�;f�$r��&�1���/���|;�!eI�O��[���p�)��+�yv����x7<��a�')�(�P%@S�8YT�WJ*��U����q�� ��Vl��$@�t����8O2�U9�|e��ō�����8S�өpQmL�e�b|�&�W��c�Vr���`�^��TdCA%��29��Ժ����_���0H=XV�U�Xw�6uI�$��>z�M��E������0`w����Z��0>�6<�O��T8�b1��f��;Fl�)ħy���u��i��z��]]�"~���+�ݿ��v�.P�����}�c�ew3S�_��a~⯺tc�0��U�ql$���ݭ�)v���K ��v���v���M�v�p�=-L�W�&CS�R��v�v�G���h3��!3�cz`���XAw,+2�Aڞ�v$?�FB��y�m�����,�ep���{3e����Uh�d5�/�F\��踘;T;P��녓�LI}�.i����1V��hG�2`��ͱ�(hRƌ��0N�3�ҷ�o*lBe�ĳ~��������|�2q:��Ē�}�?��`UF������.@��9�yPp��&"b͍��U]��{�/p$M:�	��n=k�;�W�X �C�I�l��Q�w�V�
�*��N�a���&�l��r���5
�-�ǭk���_�0�u�]C^tb70���P����h���K)��4���H,<�2­�%4��J"3�^{����,5����8�d��dۇ��i�����`�Y��$��p�K��9i�#�P�0o�� ��i~�� �I�ʚ�\�e��	�Ġ����z��!7���Zԛ���Ќ傂��DT~�.`gF�1bV%�GG?�@fz��w:���7��&ǿ
�6�x��:��������|�҄����R;�o\�*����V�N
����=�wP�S�������
�$��Ҧ���(^,x޻ܿrё��|�b	�ݣ��T:lp�M��^�?�`�W�������S���p0Pa�R�iw�K�)~�I�3qڸ��c�Ԩ(on�u�����3=/|Q_�����:�gcS]���9+7�k�/�N��k�x��$.�9��#e]�z�"��ŶC�ڽ�B̀'e���lk�?t�1Mq)g��5�@�=B�+�*�3�_��T��g�A�v^�47�"u*�GG|�_���E�(�͚D)�� ��O�e��Bva��KB~(�}V��D��/f |�u�j�g6ecu�F��Pd��w:-��a-��W:���cf���:Xp���mr��y�@F������{q'j}v;	��S�T}�aH�T�F��Ħ?�o���aq'�����\ �i�-Q>;�i�룸�H�IJ��Q<�]����h�T�C(���b<{ŀCH��C����" ��s2;[��	����h�5Ƶ`�jMV��/m�`��wk,9A�)m��-1r�*ms!�_�i
M��vڙ��Ƙ
�/ss���X%i�< ����S�h���a��A���3M��+�1/�z!�ì�}�I����Vu�ң�b�~���m���q�*��i7ݣ9A��х��V��ֵ(�9�c>�o6��(�:2� ��ڰ�UJ�升a��M�=)�|�GzFbfIΟ# N�߆)�A3������Ix9LZ��bU�C�ڂ����і/+x_P��p�"�c�O>y��JN[��-�Z�y�z� y#�S,	�k�2�^�Z�˥�撤�3�Q�1B���CĞ}�c����{3���)���t����Ag$�R�S2��8a���U�ΙSZ���O4��ņ����B�n��@��;p2'w[���â�hJU�a%���:_L(�P�"���\��h&�a�}�Z�!}��ܱ[��g�$o8:<��Z��(,��'���j��$������	R��-�ʚçU�=�*�;hyHD�^��I��Z��Pt�,W�Mp��>���/�2�W�'�7�׏�`���R6��Lx��� 
����]�|Ǔ메��Q,� ��S�}���w~Ͱ�;_�{�)O�8893����&�I��ɇ#@�,�g2pmX�U%��]:D0��
��4����iv�&����
Uc��=�_)Z�X�Iw6 �n�&{1�2�kW�v]9Ɲ�e꽥�L.8�B�^�Fe���!��Y�|�D�fl�]"�Z�����C�����Z�4��,�ҩ;k�ձj�ᐙW�F���btbն��t*5�\���K 3Z��t9���p��Yq���� ��<4�p�N��֠읥���
G����#*����85����i�2ˈ���E�k|�5{?�?$�-�^/�N+O���}DD�� ���/�`Z��$��|���۟p�گ1�
Tf"�N����	x�4J.�����m�G�%�E��u�f.=Z��tW���~�uH�
=�!6渷nt2YRsmܙ��¨�U�Ň�x��4���L������rcX�:�ؕ��@�$:�kL���F��3�&���I�"�s6��A2�����9̡�=)_yF��#��~no�3��.��2Ú��)27&hZNtp��B��>lK:��se����d;����Sг0u�<��%0� tN!��x9M+8�&��/��k�8�����~�����c�'0���7�����2p,U�y��h��+@�wg�B������v��(&yHkc"��{a2�ݛ*��������	����,:t��C�j���k����(L��!���pp9]&C�#�&�X��	�F5��7�#7
�Gr� �G�4&6X%��������WE�@�r����N}�G��}O$Ù�%|�g�0�%,��zG��hO�}�{�d�M�Z�t���69���p��+o��uz�d i}P�O��J�����D����
��ɮ�D/}��8�=���xQ�!-<Ӆ�����S��i�F(����E��Y���)<�P6�&q��eC���,y�f�����	��T���1X�x���%s샶B%6�ڣӜ�u9I>h�N(Щ�
wQ��3�Q̻_��Y�J�?�AO~����:�R��`�B��]�r&�%BܢO��0n5�����#Z�4�ej��KF���}��
Ļ���G������,I�u�\�+�}S�͌0Xn@��� ��a���OpԻRj�9+�h%�Z#���{z��Ә��tWN��A�j�\��Ői�pt(N�� ܲ�3�/�h�|� �2Ljdat���:xGEn�b0�L�j����6`���N�2X�o����:=/��ċ<G�������6pO?/�Ǌg�~\�t�&A�	��}ܜ��j���0�+=�J��l��<	{Գ�j�=��n���R�̕�7����u.=ք��L�s�ZĳK���/��yN�d��|��-��%�)�~Z2иmvO�Kw���2VÚZ_a�3Q٧�
��N~���C���_ӗ�CR�\e�����f@�l�b�
��R�}�cD����z;5�*a��N��U���.c��;�	S�ا�r��gD1�@x��J9��
�3�ys��*5�Z����4�@ϵ(WH �%��n�)%�	�V����Z%� FYT��hy�zf��^&��������_}�Xۊ����5��5�T�Fx���H��g�b,����%OJ	s8f ��"�FJO�����!��xT�uP�v/$C�R(%�Ohe�&������nZ�����}���Z��*f�T�E��n�Vu���َl�K0
���&��+|� n��ηuv�nWJZI��Q��^���TYt&��>��ȓ�Z�_#9m���lb|qɮ�s��G|��֊38�����HT⦷]]�K�8�%ZtИ:��b��,��<��R��%T�����Kg�;ޚD2���t�DM�\O�N]�:�S����iz{3��񩉑6,�Ϋ�sDi*�ذ��'����5�Ip"�T��*	�=H^ M)�l[�%��p�*�!�B�X"�X�=Y�-�R��a���|}�J7p���:_�{�����u���n��C������*B��m� �O�z��Or�'���6�m�����ݼ�eɯEՒ�_���i��_�A�I�;����,���� -���*{��W3�9�O8�H��ZSbCo����-.����M#5Ik��T���uo߆_�ē�yv��2©M�ݝ���|w8/��2�����?z	2�bXz�nA{��i�C��J�;�� �
R:nF�?�]��UN�\�\BJ�R�	��o��\y�٨���#{��EDm��b�.�U�˓a�l�.�H�x�`*�f�u�W��3�z���Gył��չ��[�{�
_�&e�0VsQ@�����I�l�T%�__t��Gm�����hf2�O�ٻ=��B�-h���/�W�C9��"��,j �Cs��q�ɭw�9!|�Cp ���8lW�O/~m�;�'D��H�*�I#��I�#'�S���Eq��Cp<�Ֆ`�Ǆ p-_��	?/�� !��8(프 āH)�4��G+���ZE�F@��𖈏����V.o��!K$���!_�\���Bib����	�@VRd~� G5_
��c�&'���U�}O��L��W`J[�a.�x>lDH�����1"O��\���iƥ;a�*�f����D�g<�qqL�k�*$���,�n�!���uw�����|H����=�^�`������ �e���u��a����)��H<6Q��S9Q�2�}�:�/I~���x���.>6�����iq�e�/N�1?j_p�7�y)` V���w4z3F��Z
�\���C5׹dI<b�����:{v0��������p�l>���x��I�����,ؑ-YiJu�b�}�	7 ��O�x �9nu�µ��@�#IkO�ɷ�6�\l�5݌P�W�C�ɤj��*q$ƎE�[^Mm������S��	�v���@h��8{H-|s8�|=|HPY�4�Z2'�فyv9��b��f�����~K��*r�(��%��� �<�U�k��D�ABDc��@�M�X�rv�����fo��Wt�G�7���t��g��#薜E?�ykr���Z�H5�� `O�[�t��#7��v9���0���Ȁ����@�)��2��h��i0����(V������B��Rԣ�#� x�A�hl���ܧ`��`ϼ�}=���\�W����.��J��g�6DH�X���(�d�F�,<��3�-(A�Rn��~�u!��5���I��h�=IQo<+�,��Y��qtk�dQ��Η���IҬT$���E����u�M�F��-&_�p ���8礸�����t��Zv�{�����L�/zy�&E���bbJE[�m������I��5���|"'�и�	�Y.����	�P���&`�F��ބל��
vs�^:5�#���UX��!i�x<�Րǹ;W:1�qS��ƪ�O;�5��g�,79W�>
s�c�^�X�A-=��@Zق���!nC�!��0�8����L*f1�M-�}����&�p�g��t�#iИ�{�d�����
�kU�΂�nJGy�e�zJJx�RŇz��B<S5��^�_p�@d�3��i_���A#}[gU�u���#ߏ�����y���;F��`�����G�>�
��2�򸢄7a�y�?v{�b3d%0�Hk�Y�-�y��;`��=Jm$s߻�K�53���/<�t��:9ȊQ���1d�Tͭ�M̈́X��+������c���z+&_A��c^7G�ʽ���?S�23j5V�>��{X8|�������*#,~�tq`L��b�;�)�xGY�_�p�mr��^8l~-m�v�h��z�p����aV���?C�k��&���TOc&����kg��ۮ�'�.	◃�a�[�8�(x.��1�K�<������ �ɨ��j���������?����������,�o�˚�V�?�#ߖ������O�Gq���_�[�OVe�c�?�<���b��0��)�[��)e�[c�k��6��'ظR�a�M���3A_��.x��k3��ʆ�\��L=��/n��&�ea��nH��@�dC7S��djc�?��1\R�o|3��wn�u��	T�H6�o��k��8L��a�����\��:���h��z/��R�je�Om���zBO�Gd��J� ��T��N�$�Av�tQho܋\:J����.�8U:���tj%w��p�(̊�jLK���s��n��@%b��
����;��!��6�1������,�O��G5�ﯔi�v�<X�t��zT�&�A�Y����VOd+-v+n�,3P�v��GS��(��vֺ/g�~��:q����UIl'Z9���M�3���K1Wx�8�T�5�P��������E>e��Y'tب�@����/�c&�=����(�҄�]���$]u��䧟;��NHӮ��nR���?p�ar�s0���/�t�c:�ƚ?��o�.&�Ų� 8�Z�5#?��h���9y�R̔֔t�Dp���X�p���1��&��to�u��I���e�%���}���ԁ4��_6�ߋB1�}��K`�ʪM���
;HVT��\h!�ɉ�x��f�����u(� ��L�����i�dx�ǆTd�ߝ�s�^�ǄB��A����GȚ&[�e����Im��fᭃ�'���ҵ ��8��FR���ܷ�����3ïo~Pgq��n����ņ�cH��"r@���k�7?]rw�|(5�p�8(~=?�z��<�3�8N�>��z "pCY� [<��Y,�ݜ�F)�(��kr�S
@��YL�R�_Hꕲ�F*0Y�~�C�J���z;��&�v�#$�j�B;��n=��>L"Uc��}�W��È�z)������7��G(}��|SE�p����z���=�'���,*��V�Ob�Y�Xj�_���!3�-��o�ͪ��H��B����f<��\(sQV�+͉�A5�,���N�/���w~�x�NJ��E@o��AX�68����M�����`�09!�7�W�ڔ�J%a/��L�*/�g�U� �y%;��|g��j��n]{Z|�!�ٯ���<&�m4�D6s�l*?��^]˔x��Xx�v�TH�h����/�j��{�Z3��� |�n%�D+9f��CaD#���ݦV��Hg��ܘ"�$�fTr��$0��y�}�A�͎�G�
D�t�ib��=���}X^w�������zu:.(ޒ{X��ib�B��a~^��e� ��G���*x}�a|��Í�9h8�aq���С�
�s�э��I�t䄹�u�q� !�f	x7��lƱ3ד���+��[ �&?����=�5���U�io�*����j��4�����,���y��v���Ɋq�Vf1;3Q�#�鼭�u�.W���?�)����@/Zn�xJk7���H��L�px��A��C�;_����Q�d	G�l�N�����>Y=�2O!"�eY8��ib0C0�I,G���d�9`;����uq��ze9O���CS��������BM�_)�-�8^b��j^(��؜V�M���s㼍�/��&g��8�KoZ���{\���.�V���k�f��JoZJ*ϋ�/��J���^`$v�Vx�;��r����i���qe~�xt@KQB0�W:v@�@<�NG.�F���L �#�(��.{�Q+5R3�ϖ��Ҥ�[h5cF���1���+d0�\�=���,��'U�
�����9��e�����V��f�)D�F�EG+�0-͛Na�a�<��"��|�Wn[(��6�{���7#;��h��^u�]~&@?7����I�3�{M�^�US�Z��$txf��4ø/�������mxas�zGB�y(�����͜ݤ%��3����`�0W��P�=]W���ۋiº���
�)t��$���̈��s,�/��a!HQIgtAO~|���d�:�O��^)�T�]yܷ����ɱh�4oZS���Ӳ�Ά��`$�s�.��n�Tā�"�#M��ħ��L,~�����PS��/� �1�`������,�zN�6n�*�ȧ�&�4tj�cG�I�RR,U��q<)QR@g��~�w���Ѐ<�ꀣ[cp���u�$�.@5���}������<����Z1��d$�A*��LDyV�.��붴:��������Ư��tC���W���xQ'���`g҇3��E�tI�ɽ~ڪ�*ߵAIh�e]�F#.+R2}md�"R�/i 0CIp�Z�i_KE�1�o��~T��O�����k7OViޞ^:��f�3�����!�r	����G� �@cȇ�%S�`a�e������/SO�@�gw_},�t���#�ď
6߷	�c�U}E�Ew�'�Ae9����]����^;�)+���K���t�Y��D,�I�o��1U��
@���;��B�^��oJ�YS�^Y1�="j����p�1(��b(c��,�_��@ �k��D��O������\�}r��<��6�<�[��̣��$�cN'x���:ør�,_�r������jXd� _�&���g����*����EYX�yQn��#8gHɷ���t 7�Y,��� ���拓8yt2^O?Ei����	C�mJ�Q$���\t�Չ��·r�����>ͫfC; 3��.zȈ^�Iگ�U_�*�Pf3�h*�!��-�M��Q!�#f��|�\��f o:�8����,n�p�<��$�=º��p��YU= �D `�m]9]K{�4��Aga9����d/���d��eAr��UP�U��P6Ɉ[�}��Tu�V��f|�w���MWp������^7�O /PM��JZ^�/bӞ�������q����P����uL!2M�'cj����i|�İ�NQ��W����Ȼ���
)�I`I/�:ܫBr��F�x	�"���Z0�5!�6a�b83 *��ŬI����:	%�/��+���
����'d���E}�I'V�&�i8].�K�旑Zǯ �0� �j]>����0F�W����c�@�z	���2��0%� Z��lEW�+�,�ݡ:�T��A8��3ltVӤ+�7��o#�����h�w<k(�s>����v�$P�	F������M�FG*���q`��)(	���E�L�F����b@~�aP]J�98�4����í&t�kg5���'�闫ϼ��J��3b  蘪��`���=�����X��?��GRե[<t+wi�E�U������|�¹�{��C���-�һ�V��Ax��UF:P�H��c���I��)T�Q��8��0H�o��&�K����B5L�F�@PF9�xg��\��+0�2m��K��V:<7�px0:֝�{�)ESpl�ce���,���N=���X����X��S�fTpSSns�*�����_�"
���n�[}jeL�5&+qo+u6��ck�׬w��L��$�Nx�8q,������@wr+��C6����Eбy��
���j!�2G�U�p���X���7+bV��C���}����?؁�H��@2M�_��X�%�O�N��W�r����_u~DS5�Ϋ<��~��_XɄ�J��z4l�d���nw��ح��N#����ם�l	�(�(�.yAE�;�t+"-^o�AK<�a?'������,O����1�cB�Z>�'��:j�+�����7��K�	Do��`f����,�12\cT�@ev^��͆}pMN*uDB���~:�;?�尰oZ�r�����F0HC�dݑ׃R�
m,�Ѳ[T`n&�hΣ�ǭ�n�ϡ�������� �E��8�'���󅭸����h��Dry���G����	�e!x�~�$��P�(��J����*PÑ�%�ں;��~T �r7b�]�}���۳����W}j#(�Z�<�8����R�6V�ƻ���ȵ"N���mIǍB]l!pxG�Z�F���6Y���X���ӈn�������Cp@N����ؿ��HR����������.eG�Z	cV����R?#�܅�㊵�qD[�=����9hgK[��aQ�꒏Z;�	J��v�̭��j!@����?����za�!����j��q�}%M�e��P�n�4��AM�!��7Fp�������ȣi4zA{���Ik.ۅ��% ����
-}�#���[=�Yk99�@M��Z��t&F���l��[�sϿ�K 	l�Lم~����|����b�r����.����nKT][��7�:SYgA�Zh�t'��������סw���p&$��
�f��^�}h&�ӜY����%�
�����s�qX�Zt^�H��=�s��c�ؘ̂�Zʔ �y��л�-E��.�*��~����7�����X��yŮ�Ԃ�;�=d�~4��`�����h���+}������N�.����ox~%�<65k�X	�d�aw�%r0[J�t�;�D�'͊#ϔ�
��9�*�gcKf�ZSc�|���9��5;
�d�NRMvF��
�Z��q�N�<�o�o�*G���H��VN���ݚ|��!�^���'7F�2PJi��R�ҭ�iQ��}�J�]��-@|]����P��Y�<j~y��&��N�u2&�ɮ?s�b�-��J��]��f�֓�yn��b���߲�@ǹ���B7z��3������>N�����`�5��Q����_!�B�R���^���8�~gcQ�2�]S���"��LS~0>0�f4�#k�R��߂��,M�|U�'.#eCP)���U�����AXy�L�{ҭ��N�ή&_9��Έ
F5ݛ�91P���p��H�༫��}�;��;A��zj�j�+�ۏI'&�Ng<����eT��J-���2N��Yp"�W�<1���T����ާa��G!�c��""L�F��x�34�͵x�3�,E�X�S�y_w?n<r�
q@���Tވh���Yru�>� J����x���s�6�����Z���Gܦn��"B����f��<�R1�b��ʚ��?�=�C����Ɨ�M8���e����\=��':Vf�Lt�����xVb��� �|��&?�5x��1V-���b�*�x��W��S��ߌb"H3&��� ��9�u
���XJ��8u��,��qR�΍ۥA�S����P���6�?��5�
;���#6�'! �xrO��v�Xǧ�$�����q�js��;�ݐ�%�̌�/��e�@�`$UP�F��e`��wݿ�m�U*���
q�6��b�@��arAU�%���IM�������t�<򛘻�7��(��ag�>� 0�Mad��kL��3υ��+h�6�Gh`����*S<�-vA���|�R(���C��z8�"U��� y�O��
����!K�@�rk�����o��K��_؅�	X��oe+� �� ]/.��쪢�W&��~�9#���4���tg�`�s�Z��[����O�؋�K̕�����hҮ��9���_�c������%����N�>�d���Ƌ4W�$eb�&�sW������jI^��L� $q��Q)�{�\1�!=����;p�]'�����f�b�
�R�j��h�%rH��Wur�9�MB�C��vH����ғ���o���%�����8�΁�F�3ꋷ�W��b|S��M#d
{S�2���M���@��N�h��r�E����_�ܷ�
�y�#$Q����s����<FG��0]����H���Ò�qL�o�#�Fv��IL�Ϸo����$%T]Ӟ��H�'�>�h���[�_�+������YiQ�D��g:`�u��RR�Y�śp�ݍ&B9c��� x��)�qs�~#������<��ik9j�G�R�V�4�:vgGmU=^���I�=�[Nb �`�E6���ǖ&c���s�!�ձ�3��Ĝ�3W�9�S�,+�8�vz�X'�xz|��/����Ϩ��@q!�15!�Q	Ԗ�貑0����7���f^j���B0W�y��`H&n��3A��ӻ/��$/A'c p�L������9:�R��o�u�������2�#&nސp��~�!e�����l�19^��@k�d]3-(XQٱr�Kx#���[�i��̮a��^�,��DU
�k-����fr��"֓����߆��k/�u�~�=����m)��P�Z~𡾶�?� )��Gdvy�O����y���)�o�X*�Ks����' Cץȣ��{�O��J.yl]M-�zqd0aޙT��8Z�c)R�k])Q�a-$����M�2
6���K��s䇞��
�T��e�q.uF�+�� P����̣J�~I��= �!�\���'�(Q��OWe�[^�������i��nۈJ��ZջQ�P�B�;��&�bP��k�^%� �$�H�(]�_]�] ��<1a����BG��őxڻ(Y�k�j�\8�$)��(�7���+�����ɱ���L���VW���:UM���e@�f��+�L������dp�Z�m�t�=@�;34)��TB�)��Ir_,0^���J�����]�~�]k!1��j�sa1i[�_���Xp\��H	}^L�X��ۭ�-��}x�
��6_K10�Eޔ��#N�p��L���p��$� `T�a��x�_�Qǭɧ��-��$������QC�0d��y��,$>�Ք=�w�7�x�$��+���3�\|���ΡQ��.D�a��?m�3�<�� �v=�e��/]��UXAɯ���
�ӭ�uׁt� `����>�R����#ļ�Ό�~䋢���_�����(�ɋ~�����D5|Ka�cCZ�� ��x23�h�5^� U�s��=��A��JϾ��YZ���Y�D��:��GdN�q�KL*y�� �^'<]8@�G\n��Z�
�R����j�c�1�>�/bX�y�R�)orڠ�đ��b8�9KQN�h{��r�L/�4�����y[D^K�Z�{e}�]5{�\ަ8�M��Q8@:�H�S�������]'�-BzCe��s׍��AS��rGp�sK��,]c��#U����e��ev�Lg|�I��֏��?경���8�m4�H�s���M������$����������	�`,� �4�lO0yD��͗+i+��ĥ_h��	u���`��gT��2=���Y��d��"���w�7���M���M
���>����B��8��O:f@{�[�5��艳�``��d��':��%�i~�c-���Z%�N3HN�Z4�[��L �8<K<&g��[,=���7�<yH�n4�O�NW6�|�	l}�$buCn�*_w��;�}�Z7ߴ�KD�[k�hfE�)�����s���lN^��-�y���S��rE��N-���@�7���p=��ɶ�x�v��X�'Ӌp����	(�.��l�:�-׸���
�N�_�.��B�MC�c��j8%���	��v��_	�y�i�p�K.cTGu�3�i%7i��e�H1�8Wٺzp	��w��S��~�@���}-!���Mܯ�
�bF�A@�*�Wy#m^�/ނ��O�'���Ul��:t�w���tzg�zc%N�f:�ꊣ�y���rU}�����i}�7�5Qx����!�as�	Cn����hh��؆�ʎ�Z0����J�^�cT땫�;�ֱ2���хsWWh0j�֛�(�ᕽ;\q,_/�緸��s��Yz0v*mڢ�܏��J��M W�ѷ}�ZV���&�Oʡ��t'm�2�DNF�j���R���3�{��F�b�}������,�p���i��ֶ���m��#��؇J�F��������\��}J�؁$\`������ ��7&{�_G��$���Q:�o��o?�y|U�|�����\PU���%�R~��]x�����n94;�X�jr��������I-��z�"q4�y��C�Z-�Y\k�	��� 9�I{#)�]�j<L{�uFU�G�hWe9q��!Xx8r(;%���1V�Hqϻ�s�F��ߋޜ7�v���Uɻ���s$�E�B��ۈ9��J0瓟��(�$�N��p��0������#V��Q��HM�k���851�4�5�( N��R��A��R�k��Q�"H�lux}�G�e�rAseh��:y!��d3�VZX�H�+�ӌ^9�5�a�a������h%
����Åo�[���#�"Vr�[��o�D-=-�m*x� ��V{��M��'l���_w�HL_䥃��H���[���i���O�j5���7Ow�Onfr_a7"�ͼW���H���3{Jz2Ja���NA�E6�,���1�r��x?���e���rqA�������)3#Z5:��쯋�����6ׄz6��2H�'��� 
�pb��?� �fx��$\>&kDY[!��iP/�:7����I&�kK��r*t���u���ּ���7��Ǆ� ���]nu]`-�]�ba����X�����&���k���p)�,�*��Ld�&�6�����uFWF2Ş6񃨫���/�Y^�Y�t&$�	�T��Ԓ�d�u&E�~���$��~�����5��s>���[���(f��P�;	~iI�W��wD����.���q27E?��u����j�FD�u�"�Տ��}az�hy�5��#e�~�|�f����c��[��nYT�q��g�8����q��k���C���/��bcmx��K=IsP�ΘfO?H��]Ͽ��jD�y�֠l[��ˆ8�l�"��38�"2�<� �1lx��5o`��q64�뎕�� V��*��<�:��|�i}?苨��cjEo�2�ĆP��zĮ�a�v�}
7.>�eڎ����/�I�;j\�5�0���Aa��d�E�Җ֢m�ٸ+�Z��`/M��t,o��3�c�a���?$o��:^��*�(y�t�F��>c�v���!�k������i�|�\���>���ȴg�?�c6��m_7���&��K����S%�0%6Te�t�����D���%Ѧ�N;��0�IB��uN���zb�7�V^�;2/ON�4U�o�@&{>\�1���i���i+Y���)Iu/��L��erj��s��cCY�I���.��{xz���z#}��b�	��0�w����zk��G�{B�>7�NB�$P�ܨ�l	�U����V���
����D�`�t�s!����i����8?2�1�`�KYk�e����p�%S���v��%�k銪t4�Uv��l�/��^���'���S�9��
b+��hҔ�tw^v�����~P�Sr��� ͤn�c�Y6��D��/tC��^��1f�O#�B<'��]pk_T�S'���1�CdT���2c�c����g���~E޲��+���&�]��2�GD�� �2viwl�N�8���:�\�D5��(-c��y�KH�]b��(�2�ƣ̕k�!Ĝ��$�6sA�n�Hsq�t��e���@:ը�T�>O"҇@�꺜8��ed4,�V%t�L>�5rƎU�Uʵ�:I���".�ls�7f�W��S95��⿪��4��!�~��n��u�M�0����h��^�&����F����p��2h0�H����,LˈL*"1�R�K�#8�����5�K��$M.��Q��M{��'v4os���3}�N��R ÷n�C�e���}�a'>-�����������o˒�[2��u�I�n���2Nm����e�����}�Z����c��e�A�p@�]�;FG���G0=�r:�z�|��_ޗf��}SN��l����+*tc�c��װF UՎ(��0i�[U'	��
_�C�X���2ud�Z�Ut<�6,����S��5�)�H3-F���a-�K�M1�MEx`�Ea��lE�Q��f���x+��!�T4�^�������!��A)-"\���C��6�ҾxX|,<u
#�*Jʽ�tw0\���i]cN��J��&�R��.��~�o��l%
 K��2�7��˼�cn�&�Pn�:�(B�9ps7o�3 YʹJ罡<���ew�4�}O�8m��H���JE&��gB��v|U�S)�F=��l8�'x��ڦ�gHSw;�榲�~� &�X���1����F��[�/�Fd�*.O/����y3鯚pȪTZ׫�,E3��`U2#�݇�Hl�y��T�ǖ�����"���쿠< k�H��۸�7��OudxK�<4�N7��=�iٓ!��}��Y�q5��eo��,�vd�8 ~�����#�>W��SK�o>�p�ҡ�b| .g9�z7t��տ�����HG׀d�S�|���-m�,������|
�rZd�}U糫_?����=��,�����!���`�0��cv�d;9�l�k�}w�r����$�����61k�������z�6��{���o5�� ��}y�H[��R^���&V��w�/���wD:�5�C��YZ��7"����s�d_�@�������<��.u�^!1O9y[j����Й�Ru��A߶�X<�m�F܁�26�4��&�CY����<x�����zlQ%�6fn�����В��lF��x!\���`���&)N!N�ap_��1>ߥP�yf��vZo:<���qNkgVFY �٭6�,t���	�>H/���ո�#���M�-�������g�})��?%WBMᕉ-�e�_�U^4�h��]���~�_\�b�3���+�U��_>�P��m+橓$���r�O��?�^n�)��k�_����όE�޿�H�ǈ���h�X�l��8$��t��^�:�/��^�
^̭t��R�a,Zo��4c�cq����&�gy��Yd+xn�C��v-!�|���Ntz�@��÷��V���y�w���vq�(����bN0]�i�s�	c�����r��G�S�HW�P���[��P���}� ��:��a�~
"ԁ}k]�w����K�oeҳ=Ƶ�@�ƈ�6c��.I�iI�O-m��z������wE��.�/��1v��׻12S�9�ȯ-��X�ĸȶT�M�)�}q?O t��3�R`"�Go�-�e��]�=v���uz!��Ѭ�M�+RIE��"P��m,&4� e�LaWԇ���w��s��G�w�!�-p�%������^�{�_��3�m�l�E�c���;�k���-�&�b4�k��7ͫ�g��o>��%p�C�:	������[\0�/�16�����h�-	��p�І:*Di­,=�Ri��!������a�i3V�ysu�im�űj?��x��M�SP�*�0�p���.!��ơ�)�E��]����F�=�jȦb�\�C\p���f*S��I�h��J�[E���	DoaiO��h�?��I?���	��a�o@��O|"`�-�D鱍K�0w	A>�j��'o��!������n�d�S�"���H�]m�5��~���_������<��[��[��%܄���I�mw����I��Ўz3����^iJY L/c�5�����k�y95A2f�'��<�b�6`V͐8��DӍ{p���C�7��{�����:_����i�us�n�h
��y�|n˳�q�B�=�(�P�_(һ9`~�`��Q13xW=-�!�t����K-��n�>Y�����|��?ݻ���lL���	���l�j�
��;�#g�@�t��\�l-���'�`K8��-�;jT�v�)�x{ =��x�W3cM3��� �{z?������ޓFȹ��!ث1u/�PI*���w�zv}�'�E=�A�;t(����L��V�5��M*`���1��큪������Lm�w�7/�m��,��&��{�Z$���q��?�'`X���Rg=�g��Q�z�>�����',��n�*���9X�U�zP��$`'�L釽Iɸ��(5�I�g�YmGݫ:VY���	���dm_�&�w6r�dHXٸ2W6��¼B�2S�osG��%�j��b]�;��5�X��7��P � :ύD�&�M���l�+s���E�K�+�Eq���-�/:E��L�3f�~=O�g%
���'�I,�������f�w���r�t5��.CQ��Lu� �1�r����ӯ�;�.�M�d��(SnM3�=��hZy�����!�����7
ɳ����5(��p��Y��.�۽��5^? #�'ґ�c[�J �J������"�'A�GO���y]ɓ>��չ�]�XZ�?(Q�^l*sF@�1�I��&y�t3��1�	]߭eV���/G���0� �beЕ��I�r�6X�T9uã�_@J1����E���z�X��k�#�Q����k&d�<- k�"�-�yw�2"��_,��'ޘ��D�������#�����^�ЈPr��V[̱7�}9�/qgF4Չ�F�떜�Jt� ��r�0&4鳦<�,`�}�ƺ�l����h�����<�ӆ��L���^\���!��|}��-`�a1�A7���kp�����&�,��N���fF�B��3�EJ5[�~ŝ��� ��*��(WӢ�E�5�C�G��d�/��b}��|Oq� $�p�� �=)��e0�$��C�>+ǡu�0A�A����\����r��r��z�}:9��͗j(}�g�^9�m8�SC#��J���;�ms�0�����¦���)l�4v�-j�̣��zG.M�6^D�#ɦO����1���j	�z�""���}1)�,�^r���c�'Dz��;�')#[9E�."�f�@�`���2�8$r&�9�u�2��B��s�I1�N�(3_u�f[ևJR�^sN�7�PQ�r��*yY�� ��t^�����Ƌg�3s{�U	�7ҷ�3t4�D�ȱ�5��;�4��ؤ&�<�ʕWB�4����(o2�&�)���|iB��6'DT��v��i��HJ%턓aR�)�GP�G.A��B�4�	^TR�Ul�2���t.�&]���|I���|�Wa�x�ҿ�� ��#�@[n�A_5�tjv�u��2�PDR
b"�Rٙ���F�L@@��|�*s�4c��1���g�Y �DF�N��p<p4�$H�xD���F���ý8\R3��A�'R�!�@tD١ޓ@���=,�I�uO�ͲPLs}�b�\���+5��%�����&!�xR�	ƚ�#��3+G��7`��R،�Z�#慧"��~ımE�Y�GT[��(hA�+��?7���ó��s2�o���@76!����C�B�����C|�۫�ʹT+�6��^������Ū�Ɏ�+�K6�9��(-3�E~�<5)�3��؁+��'�4b4g}j��/�T(Η��ҷ�Aݰ�=L�2��g�=�a�%tWhd��3P�h�5�oOd;@$E��C��$'l�	j+7hh���4y3`���Sw�Z=���Yi�FvJ-��!�}bj�T`�?B�@/���Jm�3���UA�̇yT�"��M��T%��p�.Ɗ��h�z�� �[zB?���&.�U[����&eN��J]Ep龓c��fJ�֞�1��m.�m*����Y�
��Z:}:���h���O��r�z	�m��P��U0d]���z��T����h*�S �Q�\~����UR��/���q�G^1�O��������]��>4_��/�+dz�hb#�V����F�{i��OtC�:t`�x��v �AQ����Y���g��HDb�'H7���u����S�k����S%V�f"Sp���1�q!_����S;��@(��D%C�f3���ѽ\Ҵ)�ΩK2V�
��. �փ{(�"P�Z�D����'�~�I�Z�[`���-$;˔�4��y��n��Ev�@��Bt(C� �BM�E6�0�;�m[��˦?���e��O����Be�9�9�
-�O����8Ϙ�!A_�@AZ��i�:��ᴙ"�4�mW�W��	�~���tlzjѹ�:�U�H�GJI���4��wt�XȬ�g)�T�RE�X��N:�Y���9�av��>�=��'?v"}���a��6xg#�����萜ۈ�]�G�5�ڒ�Z_�^��V�r�+4����D��N눓'$�d�Q&�0A���-�Ø��V����̈́)�߃��I5�n6l��n�����L��=4m%��0rrD"�	US	�vbKɶ��,��� 7��"�*^�K�&J��,G�taR�S�!D�d�u;�Kǰ�*��ļy��0�mL����jC������_�25�+w��xT�_��|���K*�z�_ֆ�{^��g��8"��g�UL�є�{ԍ�����	�B]�%.rZ�',���B2q �j���F�.'(y{I{qo����Vi�y��T��,KRɌ�OA9���&�%ȕ'Я���m�ݰbjR���_yX`��3g/� "�ꍅ":�Ű�1��۬mW+d�L��!��z%���'�r�����U���?������!z�m��؇	��bm�U}b����b��`Ĺ$�mG0+O.p�q�����N~�� �g�x�?a)����'K�(�+^�0QG%��2q�S]��<�_)���~k�>�1��Y�x���� ��<.��_&r=�A�fj�e�9�I��1�3���ƃ���:�,��n�ù��ٺ������ن�-���mO�.��=��L ĺ�W���׿}�u�7�����![j��,�/o8ŵ&�r� E/�U�����J��~���X��<H��,~�`e� ����>l*�����k^6�#��d��{,��Ip�x|fӈRm�1ΰ�م�ps
4U'@�;6�h;�4�8n�4��R�q\k,�¬��DE�Np�]�������(�ܾ!p�-��f�F�Vo���?4�y�ț�8�awfU�"^��6����`R��Z�)Fd�����S��_��L�M�cl�j�j�O���V�����R�Gp���XE�IkC�	�Y�J+^T^�r:<p�U�vz�t����4�e������1�{�:Gҕ^�6�o��)�-�o����Rt/���`��px�1�1*�*z�
�����1��#�H+Rz���TŹ=�R���6"u��{#���l�:������bO+C��L�:Ϯ�E��P^�%�Lm]��--�C{�"0C�q����1�#?�
XWF�'���hM��j�ʈ�ԧ O)F	�C������V���3�.j�ߗܿ/lO`J_�z��ξ%MN|ܠ<]W�Zu#GN5�y?�Ma~H������`�ō�N���Y
�Wc%L��a������;@�V�!B���H-�W�;��-څz��ν��(p��7h���>ܑ��t����v�H�k���O���*:��fa@vU5��T.p��1��ph����o���A�5��j���������n1��I��'����G�v��q.-ȸ{��t�9gt.��x{el�1��)���ޥ�d�l�ɍ����TF	�b2{5�$�&��̠�&M��y0t��M��-�Š�i�y���$����%���'b��#�P�2�m0NM��j���d�.0+�:�/S�|�����7�2��v�p��F�7���q�]?weff+U,�ޭ�+��,O1�M�b/�8086\�^������:���,˖�bA�$;}ۛ��� �"�N>u�q��I��񻘟LV6jAXJ0�D?�߸e8Α�J�P�y�=1�����Պ�m���3`����I�jt_D�x�K��7R��u�@&�_��9A&��C�ݦ�XX|���I/�!+z�xв|R��=c���&����[�^\�Ϊ���)��=m�$x�$�\��$3�12�B��#a��ϥ�����O(>�1D�>� Q���$'�j�tRnIƒ�IC��>�QH5ؑ���N
�G@��k-"�(E�pC�y�{3�R3�_�
���R��!az�s���y���[��-����xzP��)��?8ʚ|Vˏ�bX:������Ņ��]d���Wn=�����#O�[� 	�UC?f��"z��C}K2��\�<�U���l|G���YӖ��[;f0ʺȿnxjp�^܅0�}�t���v�ƥ���\� ��+�p~I�-�}$h����C�<�1���yV���C��P\���=�X�Ѵi��l[Qr���5�0A��{���M#�!#����&I&�d5�h~��M|�M��{?����2PZ�_DN?6z�ۖ%�?|�q��|7�C ����(.��an�p�� ��b�(��0����#0Tݜ� ?�yj���*��9�����#ޫ�e�v��@�і����7r3L|����R���;�V��k�k�z�C�����4C����e���+���F�L�ܮ�TD�A�w��Ɠ�è���č}�s\҄�[4W��'��ah��W��#v6Y��~��^��� 숬kx�g*���ܿ��UX�<��P�L}������D����~�t�q��'%�̍���hh��?V��<�P�.����Q�__f!����	$�M�j��p���A�J*���\�5Z��j�L�M�l����<�k�g���X��d3J��VM�^X�%�����R��p$m�7���m�v�~�����lL�#b�Z[�#��v�5m5,����_�/�����-ۏR����~�Ƙ�H��t�6��0�/e��q|+V�,y �������Ą3X������u��hu!�}�Q.[�|-������9��<��i�:8�����ȉ�&察������D�fВP�k]FKa���w�m4n	�?OV?p��'�����)�,�9JZ��Ɵ���T�"0�ʒӕ�[uf$<��Y��IA�քR�w��)L[���;J۠#,�ɉ�xW��w��S���A`��4��J�6�*��3>"I�9�ѳ�%��E��0����ٌѴYT)�R��n��uP2¤�"�L�a�92{�XᲤ���6U���^C����3BJ%��!;!�K��j�dG[	<7���=��8���)@_PEr1h�l�i�D���v����Rh���$8%uL@9G��&�$X�������E� ��	ی����5�Nn��|$�������<T���g��Q}�1��ǘ��L�$�����c�[���'+^��K)A�߱�8�E�P+Sz/���[i,�Ji�Iv�~�z= ^Z�]��� 4hza�OT%ď��i�Q��_G�]>�y�㽁�E��ž:*uZp�}�6��q*[\��v�pW2�Nֶ`}�J ��g�Qέ�gW#>�iK=��:e��0*
D�0�ԋ���th2,���{wG>���Jx���#M鄠Bh�)�z�R*|��Va����G �8�Z'i.���ژaS����W�R�M�Ju��t�c_����Pu�)�v��y���u���᳷/�Z�#�#���M&Z��y��pҦ�x�%4Vd]��涺s#Phϗ0�B��2��nd2�:RZFu�k@ԏ�]���v�rk��尲�/�WW]������n�B���Bv����Id4�@A����=a-�R���rǁ�J<.���<��$�>A�Y���"[i֊;�1 m J �eJp����_�o�n@����>��d�I�u�%5��@X��jȲ2VI���EJ)��� [�2A��;a�+cE����'=�G��8gJ׃�ߢ9�J���,RY�PD&є%=��f���%�s+���-�#���`�j�W�Ŷ�=+�	��d�	~��c	Hf}g�YdZ�:�T������t`E�eL	ᘺj.vyv�!��5�~���-.���I��ߍ�l9K���LJ*s�������P�Y�jC������o�O���b.5\�HkH�vo����D8�$3>*�Q`| �̷0&���v�_��_T$�G�	Wq�+q�Aۧ��^w�/%�_��(�iīO��d��R�[F���	ܱ��;H��`����Q�Z�U�Ρ��=���7���e�	d#A��7���'e��΀˧~�忒�����׊�/�p��+���6_U#�qbP^$1c�_����w�Ё�eق��:�����Sq�B�z��>���R��/n>�����a\J¡�g3���PU���xc ��K\�N_$!W�jp�����y�v�ݚ��DY$9q�4���U����q��/�� �������ќ��F��&��>��^-�l��85�;~�p�|����3y`*0����`I��@�F9 A)����%��IH�(�{��`K٧c0��Dl��:f�,N��^P1�G�\eb�q� D�S���R�
�AmBn�r�)��U�QH[���)V�!�n�M�T/���"�ݪ"1�R��,��d eu=z? 鬒�v�I��a�2�����'��W�씈��4��\�pԄ�	<M�a�.�`�v���d�{j��S**/�#��l���k~lj^�V��w���Ɗ�u_?�� �?�h�r��e������L��W����s�Yժ\��F�M�i&�#m��va��
&:��TST�����E�V��m̋�H7���ѢY�� t��4��i�:˳`�wR-� Q@��J�4x��h�~���șa'ëٞ]��OgU��ŖD\]9X/���jQ_�E��[8�T��1_k���e�m��2y��a;�Ȳ�S�+�!��&I�H9�y"9��sڮ=��/s�a�; U) ��j@����K��7bv�޿%��:���!]vx����z��~����bk�����8$?*�x��������*��zy�#�>ӐB�����Ƭ%���1�04l��ey�wm�,��Դ��.V�i���m�S�tl���O��d �H��
n���/ g/:s8e"�œ���;�9\"����)v�O-g�B�[)�*�2̉���{���]P?��b����ζ�ia/@�r�#[nt�#\s|Y������*!Ii��:.QI�S_��g+�ɱ��	��p�Y�Jҹ���FQ䙹��ن�q�������'Ӭ���N�6�:���<�tK$���4	c�O�R.
���T�u8�,!Mӏ/���㯘�h��Fd��P�r� ]��%G"��u�tFF�}�$��a#�cO�RqDw�L��4��%�q4_��x��a��gItD���T)*`|��g}��,��!Z(���8��{m��ӏ��S�O�Q{&g2�F��d�n��H/oq�6*6B�g� ���W�ҹ8�E���.�w�'3b7�����0�c�2��U[H��$a�a��ْ���R%�����<<�{��̹q/l��|΍��;�O �I�C)���ѵ�Q�3��o�L�ٚ
T�q^��-C���|"���tY��7��4 v�L]�\82�Є`�n(�cG$��h�����m��a[g>RH������2z1���a.?@�1�WҞ�N��������JG�q��
pS?r6�62T{i���h�F�ٍ���@�^I��?a2?���|vn8��\�A.�rW#d�Q2�*���h�~D�a�#����#:��ZK�IO�\uAyO��+���&*�	~��ߑ�+��5�ոچ�x<��q*z[�6�[g���۔H^��b�r�����@�xp\$A��F�o�����K Y����1v���+����g/#�4tg��z%jNں�_�{n��q:l���M��q�!�|�h�`DX�2�~�?�k8���7r��R���R�V��0}h(��u�L�ԁ��\=ֺ
�iB
k7��r����H��y���J14X1ie4���a��!�� �0.�S��?������;�b�cع�-��@���ϛ��p���Y���*{�݊$z(@���lį\�!E~�{�8K�6��Q�����|�?��S d�Di��y8�3S�P�M������O�V���"�&\2�M=d���Hz3�����k�k�B�ń���GB
*�4�Û9C�e�g˶��ù�D�XU�������␳������)�g��ݣlf83FDb���'�O@�hގ�����j7�&2xCf���ib}h�;������5Xؕ%�wۤVb�l�,��^`{s�ߪX�4w6B s��&YdC����X�����ii�#��H�F:-(�7�Ǚ�/��3�|���T9l?`p)h�;�k?�k�p���,��I�gp�@8]Gڑ��� L;���7[��EI%�yr#])��ߙ>���O����(�𛊄��Ɇ��fA�~���М������[�5�d������|��G}MD�U���c}�`��g*�k|��R1���
�k��P&sUJ�#ZDc�6�f�����'���H�E/:�+����A׹���^FL��kF9�d~�9F�[���5���"¡�ǩP��(�Zj�v7GȂ���!��E˃�W2 n.��bP��~?ZR�%����>Y�O��^��1{��`�1���G#�K�(���iM(�U��'�vm�v`�6�>ʞ������E��q[������J�F�K<p	����h��o��M��
�(�]a�M��+�)A��3O1�y�p�4��s�Ǟz������j� ^A��<C�,ε��y������/����ݴ���D��2 �[�kԝ$K�H��v=
�zd]:���{���m&%�o
F����������)!2 '(���]Ǉ_���^R7�^4J[W�}����^�k�S���<"s%5.>^p�~+�����CMg��-ń��I���=z�t��d�&�h��y�K��&���j�|�}�	��ǻy���_��ܶtq��Eͭk}��U�~G��/-�?��Tb͆h>~8/�N���U �t��*Q����Z�����A�^����Z�8Ӑ�X����}� �iw����TxM��?0��Qť��Z�˗H�5Pm/���9�G6u��j������v�֥�F�`�$P�=��N��6I�� A?�p�C���+���gXE�¸Ju?������8��1>�?3Ten�U�%��5Z�~	���n}_���[��B��6��Ͼ����9NYr{=����f^������V��恊��א�s�+���K��M���1�j��o
��D/�8k%c�Z[^q���R@��|�i���J��h��]C���r��Zy������OB��9	��G��3Y�Ӂ
f-T��4�pl���y�\�}�>O����u��:���e�B,��������q�N0Ϧr��9��4)s�Kn_]�W{�bN0�-?c\��Wj[�#�-$ �ņ
ɝc�妳/��V��eK,��[B(z�q!"1�z+����p��`����>�v���J֞�G���(w�]�W"�>�8�t�V�N�W�
�c�^��t�|���Լc?��\vJx�H����N'3=C�J�����W��@���cE 9�XA� �m���Q�RG����n��ZEa�q��ܮAc].fǾ`t�9��+�@0�L_�/�S_+U�b<�ZP�L(% L:x�ǅ.��O�6�_E����F˺����>��N|z�Ǒ��� X���7�s�φ
yT�Y惄F6X�W����AH� �[�O2��ʿYK!lp������M�|"��g��Eı�N^�=3m0f�$$+�KZ�"��g�	�MԷ�`Egs���N ���u�ʖ��������犐�����[G� �j.u 'V~us�@��HN�������)ÔV���GV�[���.��|c��>�邅6�V_��dEGd��� ��PYm��(zO��scR�!8۱�rbY��|��"�jӥ�ɷ��������F�nV�7Ô,7�6�91�z�G���j�z��]���7"�Y#<x�(��h~y����[�Ś���� �E{���5	��=�w������[�B�d!�TZ�%P�e(F�
se&�d`t�RQ OHrU�3H-�X��������)Ұ<шx��+7���ㅴ=�Z�fʥS-�#��`�nt��L@	�C����@�7���vB̾û����BK�M��ѻL��,�m���Ȣh�0D(1~zQ��U݂H+$�ǱH�%t"��
1~?-��yI5�q%�����'xE'���|�zL��ijF���T��41|���t���������mM*N|�`m�=ƄY%��nڻ�hI��ş1������\��j�r�]��+�Mx�5XV-ˍ=☫������_�=|U�1z��Vj(��zW��S���|�侕[��.r�2Χ�_��h`�@�-y���c��b��"z5�婔����>���x�����fHz�^�+�@����0*�ZEv��#[X�$[ �d�-t�cz�!ͮ����x}x���ޗ�i�;�o?��o�Q{P]�Ɓ����d|ev�}�*�׏V�0�Qǃɤ(w��Ǯ����Z56
�k�HaN����Ǫ�r�ܥ���%��2��������o���G�����e��IK�7~2����TZ�=����pP�p<����p}U�ם�HU� �����/Xq�S���Wb����SfJ�}?�b[��a&v����S�]���J��uS��㡕�D�r�ʳ����Ww����0���������^�X'<R��:;,�N�tGa��3
=W�W�H1��n��dt�8Ѐ�_�܄&����QKh����tgiCq	W�ڟ�g��^�yg #��1y:C_�{9�~C$�.�T(v{�ݶ,˔�nxW��a�Ap��<"F[� ]�5"��5D^r�ْ�z���Z�A`�iZ\SP�x����N����΢�-lRa�����p�5`{>X����e%�l�KxC����A�-�y��g���H�I�H�%H�sl/h/ �����"��!�D���A]iu?� |S/e�',	,'O��(^�]��"�l���a����s;����S�>�r��>�Z��`�t0���Й�BG���xSk��ڕ�HR�*���Z�P�����R븉H��qͮ���ꊛ�U�f�Co��F}��Ց޲{?k����f6��u`]UE���KG�E"%_D�m�U�C�{6�C $*��N*k�·������y+��4J�n=�@���&I����d���ނ�ble��hG�¢o�W���)̹����*0�N�(�^��k��J��-��P�e�φ���~h6ӹ�s��A]��)Xң�����YF��I�Bj�Č
�<׷-`H��y�]	�|z7&O����Sk�~��WD�o�(�������B5�}�����m�-!����@��_Yܣ�csrY�3�N'qP.�b�0��7C4&�L�������Za���V��@0b�Bž �򀏛"b�f�8�P-ʇ�Ճ��H�_б�lW|������L��#o��37�7V�S��?�y��+U�[o2��BD���b�=uX��$J�y�w!�wZ��K�a����Lᵊ�"��ԃ�!�(Bϯ��$+́�����;R�
1x[ wS��F*�|� �y�)���h��WG�}�-�{��ּ*���V�U�nxG���I4n�^�|�o}XЛW���iʶ2��"zK�T~�ck/ȁ�@2�P��f�.�^�2�'��7��i�â�|xk� k��^P�NG��x���OXxkײ��wߝ��ccc�$v9H�2�P�y/*��A4��:�@]�Ty��^�;�Tg4D�y 'e����::�#ԋ�	�ݻ�;����ҀU���B��.��b6��e֦�̌�KA57��iu��2/�V��F&��V��{:^�� �b���"S,��l�m�6�ނ��}���/��f�/�ޢ��5�@<T�\��o��5��Nۤ���v��|HYA�`���;��l�̝>i���e����K���}�W�U%J	ǲVSI��4����!u��h7�z;�	"�{w���~yN8��~yuٗoq���N���[��^х6�f��fL�hMS�/>�^'�J�D$�AC���~�:��*/u%+|��1
��F{ߤ��Թ��c=?�X�U���ST>�����F��vP���ѭ�l�ɏ��u�d������fS��u��w�
��2��_tL�XcC�F(٠~^�.i�ϋƔ�&��L�Oy���q_->�L�t�Cq\�#t�bٹ��q��n�9��OÈ�y�$w��H�FZ\���k�&եc�O˶��~���x��-�;��[��U7�۽<c�6"s6�.E<�#���J�
qBq����h߃��� �(���>p]��7!W��.�%���T�%˙Yj�̣��I�غ��c�����_�T&5'�;�_z�T��e����C��wI��L�1G�� �ֳ�F�洖aD��j�٪s�����j��z#"�O�a�E�e�d9��M��S��>��k��x�é��Tڕ�o��b�p8#�〦�Ǌ��'�pR�U3�kl�����$���ܹ(*Y��$�7V�$�D�]����\�ۭ��\d�,mFK.u���6�"rB"�{l$�f8c;ψpǎ�~/;��V�i�,͚s�#t���ĸ�Jz^K���ۇ�XI`�+ᢢ M ���k=M�I��9�'���K��|��M��e~7%u�@Rx�?�g):x+�ث���Q���r�EqEEz����a�������W�F�:�z_��']^�J��J���z��<����ҝ�3[%l'��1�kV)P��m;�U!=Q�v�~>��+��Y �=M�����6D�AK�(�R��f���މ2��cm�Z�I(`0��������ퟪZˠ��O���7F^��Z��1���T"�l:������zC�`�Q�ݎ|�:�q*$_�Z!�ݟA�0�U����-E(�A�-���R���kp���b �������??v�22�� �.�Q�`~n�zڝf{Wh4��n_�=p �u0�3��΀�/D�Tv�˅qW��?rB����`O�=�pA6�R��A�U�ƭA�>��~��X)���q��k rTKD}��E1B�$�����%*�T	goa=O���G���b��j����W����6�f&5h��g�3NB�����v{����gT��M
U�c0?�I��; �qx�hq�]`�N(M!�іJh�mu[N�($�C`Ed��	�C�5WĚ�ǏE��X>D?ɔGeV� qW�k[��+ع��ڰ2�d���uj��:T���%?i뗏*���@�1�Z�<���S���u�m=9�TL�u/��F �����&ppV&�����J���

l�b�$�n�Sv����dt����(�P�KF칬�@���.,�q
�Y�F��Ѫ[� �n��۠�i{�Jy#�5��<+N��_=q]�cyp��0	�FWg!�z1]�Y���B��O#��j
H�k�M��a'�d���zf�a��f#E�nd�Y��_�4ԑ<-�\�//�f"�<�J�W�N����G�]FTڿk_������d	��X<�����0u�ť��rʖ��CD�WʫJ��[��RH�8�[��z�`S�],���1˔��%_�C"�;�]�v��)pK���y0����5+d�-vq��Cw,&ӱ4����K Lޝ� R8^UL;��c^���J`�"���<Iq2�)�b'/F�܆-9���)_�gj������F*�+i�v�`{O���'r��mӗSڮ&X=p����Ė�3�8�cF�����]|l������iЫ\�S2��͝�(�7�� ���T|Uei��M��{ٵc�va�A�� ���JݡTʿ:�QA�m��<��R捋+e�c'�-�7��g�?�RI<k1} zx����Mp��ᅣ�_CΡ<)���!�!3v}��5>�|m=ו�]��f��CD�8�i)�>B5�@1���e��86'�����+��{�on����	�"`�ϼ���\�ø&��ڒ���T
ݖ(R2A�b@� x�"N��?�D��hJ��6�B�&x<�B�@DSwG*�6��ܥH�?���{`CT>G�fD���8�Y�Vm�[;���CK1~��)S#`��'��x��N abtS>]�&݀�Ӫǜ0�Uo�O���흌LS�M!~<��@ʕ� ��"I�{�ȟ�NE���X���b���z��ڽҭ��u�f�e�#��H�&bu�Qsj���jSv�q������a_�Hx-R�o�;!�\ G'3UX�D�6O��?��E���^:n�r�����bY������ܱH��sz]����_�`��:�BV1�"3Ɛϧ�?s�$"�vҴ�!$ֻ����}Q]�B���9�	�\E�	����xrٳ1G.�;ǝ�]���ܚ��
��t���x��hL[�����ֈAe��i�F��!�1$G�}�h���c`�Is�l�dL� �f�/̭����dS�\)�P�	�.v�/�ȱ���)
mU�o/#cp4c�f�?�H)��4�+�^��w�h��o�o-I�B��.2d��n8��:���Bu𚇁'O����RшS��U۾����G!8�ұ*9c��dAi��,Ty~D�dp��Y�9tpN��_a
�qw��Z�Dw
n8Bv�Z�tx�)@!�)>N&���~��uD�z�k��ű�<���j[U���xSM��q�.0�{��mtu�f��6����T.�>��*	[��mhM7�U�5F?���;���=�]m��}SD���Y��{v������O� ���.ݘ�ޓ��E7�kz�-$ITt��|Ԝݺ1�<���EV#Ӄ1�E�Æx"��u�I_0��q6f�a�x�2ݛ���Z��N��>^#.N�Z�k�z=��/,�	�Q:I[�3��q�@@K�#{1 /��[�u�L U��γ�LƄ�k|Cl��	�f!X�xV3�b��0�EԧE�ci~���*�q���2y��� u/�H�H���+a�a[��6ɝ��,�ߵ�-��Ơ�*�KX��䦋�C��u�*C�>Y"5�_?S~�Ƌ�6����<�����3�hT[�!�8����eL}�wx(����d�v�.��N]����X�~\�y7iÒ1]�M��	��cJ�/C�^�pu䊎4,X���^.V_Fd,�Y-[]j#��D�k��4�O�p}�rΤk�w�=Y_p�,��	d
�ChM7ن���8"�����*��>�TP�::�露�dG>�|����\(�uR��{Z]�N�*sU!N�m-(���?
T g#�MǺo��$�G����Q/����[��ѧgGax�
��\���ց����*V�0��ؾ� }>/�����Ck���Vx^�,��o��-�M5���r�y$�o	��cU�Ft��m�]�W�����H�b�2r��8h�D	��IK�`K��4�`%�;��tR�s����~:\��~��%6�L\;Pf�ů�4��	��}B�!���s�M���y|����H�j�1����b���0ܝm��$`͙oǨ-�q�ƃ�_u�Uk�dɿ4 ��O1�:KCO�K�7�O�B:��-�Z���J.>����P��م�n��g���c�.�ƻ,��b��������%
�D�lW�R2�[)=i,V�4^vP�1��j�O���I�R����#0�8{2Is��	���4����r["��x>�)��$�����_��	�)����h�)� � q[ѡ���^�c��45Oef�~�T��f�^}�m�`+�`����~�VKE�b�!M\�>��Z�I��~h�U���q���m��30��>��.P�H��$���>m�,Z��P���}[!;�y)�PJD*[ެ��� ��+���k#���{�!�ҩEV쑔�w�3�f�1��u���?@LĽ���cT7�����a�g"rp��M_��5qK݄7����N�jV�ە��S�h*��EE2Ǩq4q�<@X��bW�RA�H�ʀ�O	vz��35T8�A�k��"��Q�+��C��o���`��X\�t5�M�jM{�ƿJnDޟ^?jnfR��.����4z����}Դ��k��O��ᚗߍ�-���Ǖ���Y�H17���v�X��s��j�ٶ�������8SGg%#��'@�I��#bωCHHc��G��א�k��Ȭ����]�W3���ԇ� h���I�O�b��d��.�	jֶdc(�{x!w*WF4��?Kq� �bn-�Q�D%��S���AAQ�%.���PD�%#q�B<4G v!\��tqS.ڱ�-���q���O��>e{i�]�b�����U=��W�G{���"i26������mC�Jǁsv
���m$p�򂝃p\
pomk��̻|��m�����{��{Om���Ɵ��5K&{P!lls�$�4@ޘ#any�L�������wo��H���gJ�l��f�<ul�ھU�/�-,�f�	fZrC��ŀH�4�8�n*�n|�Q������G�N���HA�L��~���E��ų{�IȖ8ݠ��O1�R��� 8��7gj������($R�	�<�B��;�f��{�_=��I��y[�*c,/�D2���'0K���Xl�iT����E1�ӝ���1!��g	<�#��EV�/]�x��>J&y��q�&;ܥ�N�>��w�%��ĉv�38U��$�U�u}�Ka@�r���!���j=��YC*~8��'S��(�p왤+�B]��ɿ�F;f���D��'�V0�<c e T(�d�, -�(������S�L|*�0�D���q���~��c[*Ig�#�$V��%̱׫�@}>�F��Y|Pc:��F���8�(�S�`y���R���K�(��;�GN�MJ���{R��0��[*����;���e_�4��@��"�.o	��͓��!��S�44����[�	\�P�L���� �TWvĵʔ��p�Z����0OE�c�j�'p�^6���|�Je�\7��F�A7��1W|&�g�;�@}w���."elq.@!��(�[���%2���;y����R��@ �Ԏ[ې��RߺZ�m��[jEx��z�/��g�`��}Qy�qG��C�Ʀ�3�Q��."'_�w0�Ujhŀ����+�Nc%��N��l���򜌅��
�L��>�2�D�i>��-c�e��X�|�=%_B�z����#`}\�ؾYq�ji����@t~�e�3dC��Z��vO�Q�*P�-~Wݮ�Ǿ �9�t]M$�(5��:G��,����jo� ��]��*0�ba.�}�aY�8�w6l�[�ۤ��46��v�}x�y@�ԡI�ˀ�''���!�ܼ@}Om�ƕ:uv��4�Ϋ�S�ĵ���j�LT,q�2��_�G>�Q#$2���n� :3I��������͗;�2i=��#�����`�Mh��+�gz��{�YU�_z�51��A����y��������mjͨ,���a�AI,��f$������� M�,*�7l&[��^e_�)�f �o���]�*�ꁎ��ݍ���F���mw�����w[Ǵ�S�ژ��v>�|H���\5xI��{w��a ��G��f'H4�ON~�<���a{�f�Ŝ��c|չB�m�4����S��0t�bG�C�F�ޥ?�vu"�~�j�Z��lP��y��D��۪ �\��mkf��Vo���+J"�V�K1��!^��T��כ?��E��tYE?�W�*���������B��Bo���H�O��}�zh咽f(Nʣ��R��DSg���[�!�=o�6ٶ�T�P&�
Z/�GX��9���4�Z5N@ָ]��_��H�a?k<-�tQ!:���x�u'�*O�c�1���ʢG�;ՠ���c�l2���&|�6)(?L7a���+m,co-�KS�)�|c>x�gA���U��F�Y�*)Y^[i{���(�˶T|H�jb�3��I��fg���7�����e_�}�H�f9a!<c��K,����nc�ܬ�[��hXJH!
�
cN�]Jg�@�l,m�ԩ�k���ŀ���>	#�=��Ɗ׭BD�-���iu�0��"H��;��ߠ�fh�m�[�b5S��aNr�����S��ջ�Z(v鉋hN�%�R��k�%�{�)a�s!��]�Z�k�B]1Q���?�BR�վ;-�F��~NMޡm�^gSA�s; N�xKF_ۑ�JkQ����|xA�`"^��x���$	L�Q����6����a�B��Z�ȣ����_��{�d��,���p�g2�<$���&��M7~���e�-��J��h�
U`cED*�VHj���y�\�9E�Dq<�1e��o�0Ņ�IZ�ECY�[���̚��
,��l��%�!���o�Vk)ҳ+��rＧ<���(�E�oƵ����D+ao
�+��ô9��h�ת�d���a�s�%�(Y��L�%MZ���.��n"��@۾�w��ӽ>�,�9tv;��|m��{�0�O`��	���?X���␔
��ɡ����������^�X@�\�N�nLX��!_�J�Cۓ.���@|��f]ڄ8T��R�q$�쏲���M�W3Hh\BsK�y)�FK���*�eI�fj��WT;4���j=ʜjI��rO�|]�����%�j���*F<{�X8L�"�����q�:ܘ��)[�Fτ��~���zsE�#a�솽ǹf�i���mX�u����`�ť����	x� Z��?�F^�J�K^�p�q�\������U�<��'"���W�A.������dx���0�4���<���A�fc���I#7�Rڗ���Z8L?�������&֧@�g����$������J��IA���)��F�)� ߬������W�Q����X��C����ie&h�cG�����;|����G�t�fW���v����Pp�A~OT�߁9�f��[;rS^~J.#+���M�Q*�	N �rS��|�5q��ޘ�.!/���\��F�!Z�b�-
l'�BM������n��� o2I7l$��2ONeҔ�فz�n�=o{�Ϸ�j�Mb�X�+����W�����g遞ί�RI1<m-�3B�k�ȼ����c7r���ˑ�mi�O�,BV�5�a�w[�c��ߞ��w�e/�X�� �_I�Z=]o%0�<ʜjl����i�征�I�S�'�ry���v�Q��K��l9d�^A��#�*L�W�D��5h��9�Qݝşq�ٗF4��k����^=���K|���8�9�ڔk����+̬�ίsk��
�Ǜ+�i�ӦP�}��A�[L\9����8��e�'Yh���O�P��ZM������l��x����pW��m���OUZy�̠��= @byu;��e*����ɠjw4�Z'��HW����6C):v� �$��|I�Tc��&ȥ�޸wdHJ��@IlRa�ڸ���u��;� ����nv0\W�)�BU��X��1#m��
 ���Y�.�|Ζ��E0z!uyzSܾ�w�{%����iA����1�������]�c�Ty��P��j�ra�����+�]��ߟ�RH�7'�/�Տ��:����t�>�C��f����`���]o7>�Q�{�|�I�`�_m�g�U�1������D�����I"�͍{J �>��bb���Q��"�n1u�{��.���j=��K���	W��Nr���	T���J�l�.<U>y��l8��EhMH5a��VN��Mn��@`�:3�_h6�������� ���U�n'�~=�p([y�w�r8���;	8�̢פ��-C��nF��P�GR�h��!H47�ìW�r�9|J��/8IL�Xa�l��[x�G��:�l�Ad�?�}֗���V�5k���R�CQ}ͤ����8)�M�.��}X�/������R˪`�NQ�X��n����8�1�\���hjy�R@�eZ%˘YZ/,ᘡ�_6��(�8��#�Z�L�r� �(0��"��
;]ܢ���F���_���>Dj	�H�+�Ԩ
9�+:8�΅�cW�e�`�:z�c��-ۣ����]>��K50�g,`u��ʞvrM.`��ww��w��>)�ϫ���1jkL�j�庱�%��*1��Ύ��a��~JA����To�?�dߢiR>|d9ܤ<R�4<��4)����1�e��m ����
ג�Qp��8��{ �!Ժ5��#�R�����Ū��Ax�Yg�58a��WMaO뮡gy�d~�W��X���N;�Kb0����$�-(�s4�oq׬�Z�D(�fh���[6�P�J�꾻���^;�7�M�����k�o������l{�k��U�~�L4�=�3�{T��T�Ӭ-�_�����u��E�$۰�iv�*�˳�	��0�+)��B�k�X�a��#�5�Is��yoӆ:�y�o?�|i�ͮp�G���[j��r-�Xۭp1"��g�7�dKR��K����&����t�G4� �;�%Be�8k�G����m� �P����t~�7`��T_��C(e>s>z�/7Z�����D�@�0���GM=��Ƿ�d�+��և��_�i���N����g�/���vZ�^+mB0&X1˞�V17+W������궑��	a9rXLl���X)<MV:�50�"cO]�����uj&_ڽ��O:r"9���-�5�]g|n%:˚�mY���KF8�9�zF��,I_1��z�|[��D��	�����Z�X	�f5����d��,���k�T�>+�=�#)+��Z�d���R���I�#��τ*��N�$� *F�I�x�K�.Λ�5<����.I����X���Δ�}�حM⿠a�"fW��G^�j�Xlʣ �j>*�����ܸ�e�}�%��v,g�q��R�� ��1̈́R[�*wη�j-�ލ�Q
�v�R�� K�'�m ��t	����/��!O�O�:v�Ci�ow�$��g���~��cC�ZP#D+��@)�z� zS�����r�Pi&�2~�P��VÉ��"=���jn�ѐ|�-G�\������e�����n�} ֹ-��M�w�?W}y)���R��=�aw��?,C	aR��f�B��si�Y@ �:��U	0�R�<ŷ�(�j�*��_k�0G���>�R<u4�N�(ݮ-��)Ax���[��?[��U�%���`d�_(�٬Hyi��� R�e�)���<�5�t��3�=�!!LCq�-˝�窾� �+z�pZ�:d�q*N[G�*�F�~��t$�ZQ�:u�r�L$M��y)A`0��<BNu';�r����*�2
&̔n��α�j���G�F��gt��LD�f*���d�#�٨��d��k�Ӣ�o�L���-s�!��#M#�kO��M%�gIx��8�R��8!��t� ~��������G_�^�����XZ�x�ũ#�H�1"��F���F����LX[{����H)y��'�x8B��MT�EYx�V�	�!���*��f��&�ט�ʩabޅ��ؚǲ�s�u g\�&Ħ�&'�b<.���c��{
ԏ�$E/EZ"��m3����s����+��ow�t?�&� ɼf�D�y�p�?�]HL�Y��O�,� kgH~tS���W+ a_!�I��E[9+�K�W���7U虎��C)������[�j�Àпx���UK_��R�k+��2Եm�L5ڶ���4,���/���b�b���8D/���
�#%��o�^��4�jl��J>
�H������k0l;<���j:�UTx��U1��O"�N�4H��0�aF�ɐ_HBS��5FZ[��d��e5��PVYJ\���>�4T�X��}k���C�QU��I��p�T������s�O˵�Y��ą���Qh���V���f��c���~ِqo`�����6L.1X��J#p8�|������6�c�8�+����`�ӝ�눟��"�^�CN�%,���y�*XH�+U]S�o���"n�jR$�+=X/���4�rt�dC^FRk3�ӭ�ȼ+C��5B���x����df�e}e%�ɳ���b�h��Q��n79�b��W��,�t����\�ޱcT�HO"m'U�;�����g�8��ɱ&XLK�h�����|�����C�OF�6�2%vp�Q��V��5�$A؉��K4��A;}b��0D��'�H�3�=��V�n��g����(�'�_�ܦ�FRI���^��ǘ���结~�2���^� ;+/ �H�b���i��)�Uh����٨�j}o��I�8W����G]���3��\}�E�{9��洄�Vn�}��������:�N���*���<��I�39]G$����H���=X��]D�P��5rU��H���&
L�=�0:쀷�|��Ǆ�9��Na�KH\ u�bi��.�NV�=G��{� ����hfUYjj��L� ;�o/B�x3�3ۯ�Ƕ�A:a(-Ws��?J,�Z��FZ��#ڛ��������c�ՙ�}�r9���J�.�N�gh���żB88Ӛ}�<!�����+��3�����9#<�NV"3*��K�G����bk۬��!\��h��T�и��N_����P�,�,.�{G�������屽�L��ٽ�=�ndy�2IRwll����"�N2�Ryq����=]��m�	�Z�aϭ�}C9z���9�7�،iz�|)٧�PՐOn;�`�}ş2u�Ņ�z{�kz�0BE��1�kT+�R������r5(�Y�6N$��h�2������k(������ʥS»�'@������p�r��i-� &�B�(Z9ݕu��٠����]�c��^����&�U�z^����F���R�>m<�l��G��Zf֖�(}��|=����p��ȷ;}˖�/F4�E�1��E�� ��
�äg�|;yY5���HE�e�y�=�,�s�((|�<xIH)ޕ3^ޱ����R���^"�k�*[�٦��gdh�y�P<>�~Z���~��s�j�t*�Q͒~��C��6����ʠֆ�tX|4{.ԥb}��29������1{�D�����2��D����Gy�\!�؎{*at��HxzAzj�9?r��_�M�>}M��`�<O5�F=C:{\3z�Fv�@��	��[�p��b�N�L��T)5��G	Y�u�9I�c�;�j��xT(h$��7�R�wqy��]T���p�L'�꤈m�k�-��_�h�D��7�y��?��ۋw2���NZM��2��z�� .P���+l�tg�/?���BE�)���_G���%��1� =BcOI��%<�s���R�X/�O�RT9�k�.,o,)4�JՁ����Br�O��\��U�V��	����rW�����%_2:"L�M�Q�����I��eO.�筳"Dz8�}�ڇDƩ�~⡺��'�w���i���8o��;�^�ȝM��o!��m�� �L�Ջ������})H��ڀ���w��"��I]��)�+�ͣ�_���oy
"Ɖ7����jxh�>��8�ܤ�L Ue��p��T�\��=�_n��D�.��;��#�ղ��~�o�>�|����Y[c-R���:sD��͵��:�X��9�]��R<�Ch�xe�a���I��%b�Y�VD�5GV��� ��%���)�k��%�HS"'ijH��<�US��?;K�)�(����_@�G�R�4B
.7�������j]bO�+h���$J��Ǹ�C�N�]�C�C����$�"J�8�F�DF/���R�7�.�0F�8Ph�h��jH���:&����`'M�H;��PG�!I���P�n%�K�%|�o��4˕|h����EW�[Hhl���nvw�I�����˃sD;�Y�'��#w��/����T��ľ1��\7m�볊��g6},	��'jM"��X���T<�Hr��C�Y�]�0�����`���3�u)�`~��+H�`� wD�)R��qQܼ�O���o��/G,Tk�<)�-��$]l~He�*��sX�{�����Z��&]
�8D�o��S%��,K��j�]7�m�#�x]��Zd\C8F���h�)X����7uS�ʛ��F_������{7�я���s�O��Q�10[�iu	v�ɪ����8A����e�u���F�I���1�(I3���RP�ȿ�hq�l�Z*R�	ms-��u�0�p�p��t�� r%ʻ��-Ьb�6����T�Aj��@e$�������&��+�E<n�#ǒvF&�&hw#�qD�J=��_@=���rE9mU�e���5������^�e��y5�R'��iPX�i�g:̝�"h\���-q�Jt�{Nɲ��r�G z���ֹ�����8�)�e0�7 j����
�+9N����se��� #��������ى�M�)���5�|��P�j�.��.�& �߄���?�s0D~�Ĥ�t1H?d�������l��f�bJ��Y���&-{(@#8��a"F��2�U�	���0����A�G�����(����6���6i�g�m���O=�n�O}�(,�ހ�gF�?}I����i�_&�-��u���7R���{M{!�I �خK��}A��F��-M͝ `���T��AW�ed���_#q��n����D6̑���b{���\z����5/���EeÜ����aF��KKy��},3���	�ʰ�#����0��_#�g�@Nf���^E����!��l���k�H3���c�;�S�f=I	�!�ht،�g���I4`�C[�|��s�#58H����=+�;��2��3�6ID���
xj�=[X������Ձ����p�3�+�u��>��m��U�W���l�E~�]pCy:J����Q��E�g�)uY�{k^�v*�r�6@��U���M:��/��[��M��Ƴ2����(^~��q&X?�hoP�W��L����F��r�[v��h�*��e|񊟡pJ��q�x2��6
���� @T,�i�����hl*�]'�Be/�=�c�����j�s�!}^�GJ��D�lw:��T�5�,����2~SJ۞D҉��>C3e2��E5 1���T��	�,Y":�^�Ll�׽��D1�<;զ:��ڲ��䜻���=M�D�Ԏ��|���I����f��8?Q�
T:��O�X���� ��-�}k@ٜJ193���=WC�Go{�F�J	2���>����k�̴EF�-�����'vC,�˼���_��Gz����Q�[�$�趷d ���P�U�f���������G��8/&��@�{]�3��6����Cz�8����R���=���ߛXe���C���cb��|Ҝ��Lht��,���ZRD+���ű�7@�Og橌/�{�<䡗&�B��%�f����Ob�:���v�`f�/AZY.=i��*�W����!�{������D���3�j�Ip˃��Y��2hA��*dm1�{d�u���.?�_ �v��ܱ�X�$���#L�=���(����;m�5'���ݶ)�W�[2H԰�. ��w#��^���������� �\���t��\?Ѝ���-�v�0=H�� ��)��nE'������|����f��Y���ψ܉�mNô?�xx	���*c��Zc����;���pO�	�/v4D��9'6� �v��l�O��c��1��&ݜ��	��V��F�>&����œ�=������~�5�)Ͳ8
��sf��,�-~���E�X�U������H��]��;��PD��~Q��]�e�Y�oO���pA`�WیΈ������y<�7���t�8�ߍn��B�54�l^�����+v����p��Ǵ�U �ی��5;���'�����(��X��"i�a��������ٞ0qa�;w:�A�zi�!��)�@�a�R�%w��Gr��h�6��r�a��SG|�O�'}��)G).�$�a�a�\�њ��
0��%��۴�b�6�� �-�⧦!߅���Z���r־SS=D�=jʝvS�#ONT����w��:��	Đ��d��+�F�ap���9Fٿ)���',g607�\�)�p�HZ �=j L��EF!J d���\�6ju���K��4����hsrH�5��w��J���bn�I��M�{��Q��Wn\Lʊry��C�fXs�[�`bm/!-�s) ��8�u7^�B<�M}<� �w\$�z�G4!|ߧ1h��A�x�w��� � L��T���z�*�3RK/� �i��j3-#�ѷ���ȗ`�����'��sD�ws\��;8�O�.8�בR���P�S�=p��=/��@��8(���_4�Z�A^=�I��|�b��V����A>��}�z���h��]� ��d0̔2�vNȢ�ID���߂�Ĥ�b�N��y��wNT
����Gxf��q��'�b㘿H�9���zg��j��C0�ZF��z�@`Ud_�����.R�Dok��TS��3;���N5;�@ea�V8��_�3�S�U��&�_&+oN_xn���G�(��%HY�[kO�M����K����r38�<$wc�Tj�'�o~�KY�nS�U����Kc?��j���Ѷ�R<ƃ|�7K��G�d�%��]��+����S5�u9)���)�G�G�_l���z]�S��l�Ůw]W�
���<�]�~n��%W8d8��t��=���U:���gsSLN�T��B����G�c[��ʜ̬mi��	J��Eܘ�/?�Q#B�^�G��_-��h��jq���{��4���'���K�ulG�*m��"k���A/@᤭#���,(��C�_����� (74ʼ��P�!�(e�7��5���8[�e�	���d[��8&�b���Ʒ��?���l
lTNf�j 2]x��'a���r4Cc�B�X��z�7�M[g��Qaa}��;�+�yp�eء��Ų�!ӗ7���wI1���u7��h�|yg���X���*ޠ���x)��������1�>P�{z�x�և��S<˩����҇[`��WT�C�nB�}Զ�/v�^��w���Ӎ"����zf��1��I�wL͑�r������k��ݿ��b���<q����ҩ��:Z��na�p�!=n��i�Q��n�2���\��f~�s��f����B �h5-Lע�+/FGq,��-�4�
�e�k�[J2���Ψ����5J�Z�9��w�H'�9����$D͂�pF�3�*f$�ف�%ߩ]��v�ߠ���d��ބ�I����`�Aj��-����w�C�P{K/��k��VJM�K��-�Bc���x����1��˦��Ne��5��먮B�VG̎F; ����i�^�i:��p�⁜���&�1�
b���d�=�nE���c\z���>OXG���Tp
���q��m�ݠm��gX��|( v���70vg���CZ�����%�ͯ0��:G�
e>�$]��W�6�9WO��:0&.>g�kHK�4�ʔu��N�9�͐be�\"����E�M�4Ф�J�c�?���-�XF�^F�9c���k�0/0H�+����=�"*:M��2EDBo��5>؄v���ـ�C��R�p�or$�\��ZRf
��v��۴��!W�O�jSC���*3gd�?��[�������LB�s6��j��+��\�Tӌ0��lָ�%=Dn�$3�����������CeS�K��m=���6�#����ՉkmW�!H�,���R�xc8N��a7%~��O+.Q�(�3�Je���q!��/���I�"jWf�_� �Ye=��[\�@G]]8��;s��g�T���s�g�_$fX�� ��Z�
�a�{H��x�.ch5{�XE���� =?�R�/�9���ԺaeDdV��u"XT��5�3Y�ϻOt��z� �BF�5��$��W]����I�N��a���o�������ZU���@�<��R�*#pg�c^�Ĳr�:?2�k�D�أqG���^s��SP�a�w��ߍ#0�/��I��'3�#�b-�9?)'�c���>�!�u7��1M���ۖ�����ϦTO���9uE�6fA-P���@2�(Q/�N��LJ;e�d9J�υM����R�[�d�"W�hS���Ø�Է����#��Ć�l�=�I��<�^��c⬹�E������\�v=Ȣ�\Y�t�I#Ҹ馊���&pY�5���<��Lռ��/�'�}'���z*��:;:��tMV�e�*�yi#��F+-���� u�"��=��y{o����Is����y>�ɢf�<��d�x#d]��T.��x��P���V��?]Z"y&�(�
�͍dkD��bf��!y-r>Ő"�E�T:����م3)���EJ:y����k��о�(-�]J�PCl1NmD;`)P@���e��0b�U�%t�-���6����o���ma6tW�H��� ͓R]S�A+�K����&�}�3J9O��[->B N�n˝L�b���Tr�^�&*Y}e���pB!ȓ�P>@�^�]��]�����Av��5D����'�{���G��R������TD��݆u�l8 ����E��������Z�y-���#�wZR^��Z�!*����W���@WC�8`#��>+�p�z��{P��YLO�:�o������+M#��mE�q�`��z#�c�t��9]-+�13��ߔC���%�fo9]�q0�ͭ:_\���82�^�h��z.��t��`ﷸ>C��ں�L����[�R�8�x��=��>|�X��N\���	WI��Nԉ�]�8��#�����f
v�l���J���U��l��¨}�qC�d<���������ȹe��x rQ�&xS:��Ǟ�e�خ��x��(��`�H�t�0�lg2�M�B%ʧ����ձ]��x�=2����t���OK��H%��q��V����܋��>�S�����b���ܘ���n�����Sf��C�ڻ1�H$��ř/b���7ة�sٳ�n$��a��uuW���
𾇻g���-�]�x��S�/�����}���;ǹp�Ke�A8ቷ�%�f���N+�#6��ZRj����m�u��X�2��p�"�ɞ#��Dۋ3�@"�~ґ�3�����lw�S�S���^�Ξ������\RF�1@r�#E�O���,+\�j�;׊��]�:�� ��j8,���r��m�T�m�.��̚����u����C����U�2M�m����?���E} u�	k��c��W�|���锼F
�V����"=k��GJ�xov8K����R�P�����O�1�:`K�G�M���=��s��Zo��g���k�IQ,�x��9�Ď��b 񓿕z^�_��8���.� UN��!6�B�ܠ>��B=/D�������Y��=�b,�w�x�!E�Ϟ�r�Hvz\�l)�'��y�\���UQ�~+T���������!�3�g��-��p�U��M���E{3�˗�6O�C)�C�����P�q��Ĉ����z�o�!�B�蝏�AHu���灱�5Ӽ[�T�|��yG��U���'��La_o�1���Lp@��(�t;�㔇�}�lA#71�?��|_8s���0/��U6l{�#
ʤ�2c��4�7@�.����y/�C:Ȅ"L=�OB���j �>k�KV�����«��ڼ�����>9D]���Az�a��{DmÈ`\÷���ģ~:qB�8������v���$��M4����] *\.	Ǽx?�g�"�79gB�o���L�V�3l)k��T)~9Ox`*m������Y��X[�Ǒ���@��ґl��F�(�n��(O2���UMw<_B9(��2�l�F� m� �s���?m���ի�.���h�m�����<:�k�gRV�㉸�gq*��{����6ǆC>�쨧���i8�/��r*�������Ӳ�1X=��I���>,[���{�Ů���FsM;U�g%�
f!��J���$K��\�ձ�9"�ٚ�E�<�-^�,���&68_���ho���w,K�o��������xJ�����?Ҳ��a�L�B��ʻ����D�lo�{~|����� p��?6�~;Ȑ���+( BŎ��AĿшc����f*�a��CV����M�%A+6�TQ�� ���� |�\T�uOy�QR`�kJli�k��-��)�*Ҷ�eZ��j�XJ��j"@`K^��b�>4���(*B���}y,�ږ��m]�":~�V��������%�64֩��r��y��S��ku5���Vջ���(�NgU�(�='� Wk�ʻ6N�6�($Ջ�'j�ã�W�h7�IzSCp�F(&��!����(�Ym�9����zTo6������B&>~�tM���)�����ңtU�7]����q��b��@�J�Ż(|�p�`0<�B�;hwΠ���<�<n���?�x�r�����*C�7�NVz�m���$����vX4Jk����u�\��,[�z��Tڤ��.��ܬ����V���S��9���;2���3K����C\���T� �+I9:Z�K�!!��S[ܚ�s�~)���*/b�����8S�^y�t=^|��"�Z'����%+��ꂭ�$����is���a��߽���;�4��G�)N�]�N�� �'�m��훬�X�`LE��d�&4
P���;�Txɢ�*��h��[p���	a��@��>��+}՞V����W�s�=(����z�xQ�vi��t�Ԍ����dx��ksp`�׳���m���z�'���T7=��ݺ`���	􌩱��U��h��+ͳ�U�G�xHl��U�Ai�+9'V��m,��Ro��!�`Mt����H �qT���P�F��b}��&C�R
�a�92	հ=�a�ͧ3��}��%������H(�#���+&ſgr?���;c�������0�oa��}U����K��ѽF����_�hP�*\���#佡�$��OYDQ�:����A4�ϳ��7�p ��R�D��.F�����ъG�mA��,�7��:\��,�R@�5�"�����fȼ4�@�d�R��
T\��"�D�K�S��C�K j���~ű�@
�%��A:���a"��������'+˓��bj�� �����C��v���~�3�L۵*�/�՗:�������QM��6T�@C"�Y*NN��N�s��/ݚU),^ZfGՌ�3\n�,R�^��Z\Z�����Ў�3�M\���[�L�8�1�zEޝ��-5	=H=�U�ـ�[B�8��UT"�n�������ؖQ�B)z$��&�@U\�|�\�||�?es����qg\�-�2ʰН�5���b5��+�S+N_��UX���<L���9S-����Y�b Ԟs|tx#���W��oz�4m��E�����՛�s����B�#h��X�Wޞ���ժ���1���Z��H��>��Yn2�1��&M�@����~2����6���]��.�a:���Ju�>H� �F�#oRB�PGP敮�l�W&�ƹ����!�z�QR�V2y3�8��<e���{��Y��4G0M%vɺr�.���i�UD
�@�;�z��mm0 &��6�afdye�d�w6��)o�,� ����Qɯ~f�6]b3��g��]����$ ��\�5�XKY._�I�D���۱Tz�i �1E���<EȘg�9J� ���~�l��0Z�"z_v��X�m����M�G #=��=
,*�@Quꭴy���?��$={
��[NR�%�Rz:g\�	ޮ���7�׭�	�m����#�ñh��]f�[��B>��X�:ږ����%B���mQh�R�z^�x�l�V�x�Y����!e�yWq>�8��}�@�82�u5U�x
D ^�l~�r�I/�ЍC�k]� �⋓�������Z]�8=��=�{Uxl���Ly���Û��>c�U����]i��>e=$t�Ka�r�l}�^��͎l��#}Q^k��k|z�dAc�]�.?;��į��[o���\|�_�A�ġ����~�����l��z����f���U«��IB˱�E~�;�M��ʁȚ�A��i^ھ��$�'r4P-~Q����+�(<���J�8s���>���ȅ h�����tƑ�3�N�@R����[E~�Rց9����h�=v�տܤ'���:G�@�Y��x���F()-
�eGL�Ly�̇8| �@�hTK�֊�c�����k	��R8\�5zD�S��<,��\�1��V~)m]�e��� Rg�p�&C�nO#`|�IpOuGVꚤ�"+v�;},Ⱦ:�sSK����Nr�8��4�?q {�tB�4����ʝA�̩��5��s67��԰��O�Lӭy��[�sT�߻��j�*�|��Ϟ3�/��9������2J�5���v�?�m���E�:P:D�F�8��O��ڬ��!C?�^�VC�r��<�����,6U���._B$�����������fy�} ���^2��[��P��HW)�%�K�����lݨ���׆�qS'��\��e��	�?����9���\<ꇆ�̆����4��C�ֱ�8�h��f�����c�����
�W�#�Kf<V����>d~JY���颛����%�{�J�5�/��Ͻ�%�m����+SQ������!p3�9�Ͳ\�,�	��������B1�!H�3� �s�9�~�b���'&�Vqg6m򣨣RA�ƣB ;rQO��2r�g�~�R11��*���mB"sS�h�C�$�##������ܼo�M��#�[g������)��!ܔ!��.�V�&0�T��=����]��!�v� '3����?�O[���*4��,�Ij6����=B���W��ȑZ@�0؎ĕ���ɝ��w�F����0y�;|�"��<�c��W��똃W�M`'�&�!��/a~%x�᧽������T��@�&�|[����7��5B	(��չ���,��[�	^�G�A:�ѽ��+��<i>	�E��	1�(���/�ћ%��3�}'��K��軎^���Жٮ~�V������叻�4��@@��)�wj�*�g��!�)y�l�⊦l�g��:��OA���_%���D���
�A�nf/g������f��q���[Z��e�\�d�0�Ǽ�}�D#5�]n�1���)b���!#����[��Es�y� b�}��VZ�䎫M�&�-إ����#|���`�ŏ�	�X�݃qM|6m�)ޘo_��D�o�K}KofV���������m����k��Y���'4f}�n;�vIX����g�Aj���gU��|��1vZ"�1u������IöJ�φ�����3O�l�d�i-��}5��ڣÍ�|A���۰��@~*Πa ���c��`��x��,t����S��B(��t b<��9_[.!!z��9P�Ƅ >��=��$�>C�_o�e�ǋ2��w�uӋ����6Ww	�Q��(�$'6؂O�D�1���yl��T�G�ʤ�4�AJ�α}o'ert�$��N �G�~.����%��;���<X�/;�SM~�uy��p����g��g)�K�-%!�i+[H����a�ۓ�o��}�0�-�����S����+K��K��#\'@p�0yg�8h���:�<p� ���*��o|2���\W�ؐ���Х��P�L���M­Kc��w������1�S�!�E��t��<���{cj�D�(��Q��m����\�;�l�"f�Ȩ
UlX�I*�3����7�y�O�]@��{���&o}����3J�-��mKh�'����+mFiW8�4"��A�n]eb�]�fw��#��e�w�o܀�����SXw�B����e���G�qS?:����� O85�q�s�j���^��XC86�o�����5Y��ژ�K�ϸ	dg���r���-��=��p�=i�����^���q @�v�kSC �l⚹�t9�$R�������Yo��p1��.�rK�
�:�b�i�l�n�R�������]�6F�#� ��3J����ϑ�� C�ˡ���N".7b��4������N����ީ[ޣ[XeNs�&�Y�(�:�fQ*H��<\��9O�A�ϰ?�ᗢ�����u7M�Y[��T��s���b3�����l?�
nfO�"Lm�.QH �\s#�̥��\�$�p���81�A���y��F,����l5[�	�E�k%3��.ʣ��9E�{��t�Nڕ]:�y׺� �z�d�������I�&E[�am����`0�΀\1����C���#���E:�&���^!�ҵ#�s����W狍��JHx��}��"�{u6�a_�y[b~~Z;�})pBk�l��>�<�~���4�y����Y����yڪ@K��r6(Z�V�ً 8	>귉~�g�F�7,M��~����M�6H ��`�m(�_�����q;��x� P�$8A��ٚ<�[�ՙ�1�7#��~�k/F��~Fn����1��`�yȲ��څE(hj��`����j�jMT!e�q=Ϫh�y�<�/�B)*^���M�A���N��lJgDa�F���Q����X䓏G}�>�;�<h���ո�����\`U[�92wq������(ڨҙ@�f)��>.���R)��ޝ)���=�o�J7��MV4�^0��X����+v���8WL z�Ҵ�h������p&j�A��4h��Ij��а��{�������H����I&��@�G�ɵ��t�ЅA��.r~VoZ[X�k��"���h�'�ȸT^}���ȵ��x,�%�#�}�M�,(k�;F�k\Q�=~T����C�W邧s����S�-�U��.`�&������5P$a�S4ª�3E��Rv�T��"z2�B!���j��Ba��1���szV���P�v�鬪�r�o�����>��oy]7`ɷYg�G��/�� sr��kڮA�ۍ|}��_y5�=��܄0��7�b3��4+r�6�or5��������v�<��w;~rp�^�L�k�jN��`�S}���yqݫ�E}�!e}
���1F����y٥�:���}
-y����-|�eIU����3V���0��8n�m!�p}�t����&_��2��ba)D�dC뭩����b.�m��Dv\Q��D��ލq����d����	�����-�m.����5��M�+� �6R���Df�\b�<e�::e��>��iV?id�}��.㸨-uaTfu���>�4@p!�S��/����lV��4[���� S�쭖+��@d���af���ĒHDsS|!
74��;�����Wa��Q�qn%=���z{4�Ą2;�L�q�X��V�na��j��n�dG�~?��9܆ҭ�w�����8ƝJϕ�0��~�[X��f3����y��8���ey �%�R���%�y��8|G��d��a�ݽ�8c��:Z����2�ǻs�:���c��+��Ei�Tpl��C'=a����x�cNL�r����h�Ey�Y.����ٍ���Y��UN�b������9�k��27�ٌ��s�u�"�4t�û�
Yr�Ƹ�kS����(��N�k�w �lc�keEٸ����h�{��v`�LT�i�&�$��[�׌"}5���ʁʑ����5�.�I;��l�ǕE����š;1�Q2	/���K�?���c~�<��	�d=x>f]{�f��(�kD�f�\�5yd ]T�4�{tS�J��'�*ϡ'�?�>?��v�p��~*`��$i���ۓ�$�䄁UD���0i��nu��K::۞�M@�/�����ؒ@ ۉ�̀d���zG��F����qY�ZW�]Eǭ�8����ōJ�S���;�k?!��c�XT�Vo4W2�^�dE��/�]�����
2#������w��O�{q�7}�!�^�'���![�hǸ��Dw!���6?�r?�$<���� �Ԥ���;RM�'��r(T�ǜVz1�f�d$c�_U�Nu�T8^�ׄ���/6�=���pi�K�:p��Sh����=T�W�DGn��fu���р��Fؾ�*��y���Ү��v�T�x��N�!f�!!Kr�	rӘ�D�,�U"�o,�C%;(��i�n"	:@ض="8e�*	;��輸X�/=�kx[g�����P�f@���b
�gz
��ö�ג��^��h7!ꖗ�5L��G=� @���U	���;�++I}Z����^ﰀOu���JGo?b�j��Y��\ꡃ�j�]Յ\I0->E�� "�S��:50҉:Ə\S[�7�Ȫ��S��>Am饫	CeM�`g)[^=騑�����u�(�/������8�x�%70�m����C� �˖����Z/2_�=A`�Dq�8~#�u���3,�Z������Z�gܑ7��C����G�3n#���T�H)7�1�7��1��ͬ 6V����Rq��v���k�ȅ�Ϭ]��a�!G�1򄁡�h��A¬B�7�^q�m@�ß���찂����'!:��Ov�"&��*���������*��I���K
��9b�1Pɂ�w�y,����.'�6���#Jm�.~1��"C�
��W����zpT��+��|�`��E(��� ��E~u�#1��h��P^����,PW����(�"1~��v�ȸ��m��<�7:����3,�$�?ywS7�&�W�B�G�=S6ތ��u��`����f�yG,[[���i��ov�
�T��1j�E$$�śQ�J  ���=x�H l!K�űN��9ч��=�UWa�s�/_\���P�1�&��(U+d8�MZ0�3a�!��Y1���05O�qb6В@��y�� o�%��Ep���滚�ʺ|A��Nx)4�A#�Cl�s! �	Щs��'����8�aS���$/5)���U��N�7�.�w�&x&K+�/A�ؘ���x+t��췱�)A�����s���w��>
5xq��,"����˲��o'�l��:6���eOT{2V���7-9�1;�K��{K������j�:�tB��l�9�}��˕�7�%3�P�|EVN��ݦceG�����p\Ѕl��`�M�t������T�(B�[��D]}�㿑�͏fA��t����t�	Z����S��[�S�,Яd`�`�@ZV����ψs�^��yi��;T��
��?Ͻ��-_�ðjώ���,�Ixa}6ώO����q���3�A��n��U ~_����4��KA,�C�ڼ.�:6�-��43�#�E�MC�0�kJ��"����z��I�t�����x��B���#�����H�����;	���R��� �6i��3�:����=a͉�W��X&&^�UB�����j��������{�U�x��vC�}dA3�Q���p�D��$����K�jDK�C���xC�_ �Ce�K�:����D�N�Z����d��Ar���+��䐭�,�f�JtJ��w�I竱/7X2kR��|���E�7p�T��&����&��,�{�-+���֝�p����`�_s�"�w	 e:b��	���R��r
�?�^�c��֬�~G�$�;��~����'���LJJ�Yք.�+Fi��Kw�V���ZFӢp���
A���j�*&�~Lܪє`�L_V\Ud2T=!y�It���<���u�U��{�6��7�w��. ���.5�{��.�Sj��.	�&;��Wa+G��6
���-��Xh�oAx�zS���X�r����u7�An6N;װ��$-��3�7�9	�z���;0~ʓ������+�#�T�s�"���O(�f>����o"9��ֹ2��FQ-�b�����cL6T�=�>)Y���ʌI��V;v�$,7��4��B
��-��πswuW��[oؾ�`iU4��������,��x]��P�ƮϚw�X��q_��Q||ɩ@sG��l�};�=�,�<ª�b��}����o'!ȟ�.�r>�>%A&��.:���p����ln�:�?���$@g3wى��g����)�W����6���)�UTw�[���d�I]NK���=�o�PU�w�떼��{Db�BX���\ThӮ�8U=�/�D�G��貜+�H�d:=l��90��~� /	nOm�^�ߒW	�w�s�8gg&�q��܎�6sR�Xn7�蓚 9�^����d;�~�$ J�57�n����mE��..��s��1(w�Pk�N��_(�i��X	`���ɤކW��t
O��p}	�T�H�|2�$�yR��P����q^��7�!��Ɯ\���i��OƒY�W��:�D��Xޘ�ٕ�^+���s�<��8087� �I2k��'���-g��d�s�m�xt�I/'+�O�����3>�2o�I�΂�׷�^ŧk�`�q��e����@��Ҙ��px��!/(�ԇ!!�`��s_Q��6L�N������ۺm�YE��P׽�&KE<�{,�4P����#7 ��<)���m�q-݋��`;s�h��N]=�k����Bl��IS��1��X�;&:������K��gœyF��9�.�$��z�j������$�LA�G�����D�����}	��ŜP����\i�*��C���^�h�Uk�qHky�w�]���[�f�[TF���Ц�o�o!8|�1�nqEY�Z;������6��K(�B7&DQ@�xƚȶӿ���,�>&������4�A2CkTK�(V3į��w�%�Xy���_�N�*�Z�pӇ���U���p:{�ÔຟD;��H}Nn�R^�����������J���3��7Ș�O;���yi�r=z��O�-�1<�C"U���	|W����xn�`Zr?�8K+��ek{k�w�>�0��Q_i�׍c#ʤA�n�0���� "?����x]�пڑ�*e�����f.�C͜c��V�ף���s��s��Pe^gUy��2>�>0i�{�bV �m�NP>�x��b$<� �\ݞ��� ��-}�n�.��U�8���D�P[le�c�Z�����KG?�Skt�D��e���8F��A�۶]ƽ(g-&A^�+g�-�S��\ Zy7x�M��pK���q�ң1�ezX|s�y�g�WR ��m���ʁG_#6�^�o�q�)�l&��ur����F�^U��n9FA�*g�΀�j�x��G.:�(p������Be�a��+�)�=����g�B\]���|-m>6@ѫc�7�FmbiG�����%�S{ǵ���I}l�7f��g�'&o�w:�
g�PG_�k*�OǙ����+�q�z��8\%5nk)����"ǆE0	����*�v����ax��F��"�w��"۷@��55�<V��8�x9�ӗ��_\'�`)��-?l���R�P���\[-@-Ŀ ��p���D{-�]�y��[�h�?ޗj�!�a�1�δ��݀m_�	�ejs8ޟqO}��+n<��ñ�)G�G믷���T���Ǒ�{C`�Y#�CF��=��a�]��p�d4��,:�8�W^�X�/�0����f�ŪА�Yp�� Ջ����0�� Mf7�R�B|��l���IR�& ZW|�D��_�0�!�6%�2,�ayR�5k>7��Q�)ל��XMLD�&I��g���70@\��%�����ܟh��H,f%F�#�&�ҩ��+�7T�C@3}�(c.�c6�Vq���L�I�'�Ee��鴳�,�2��*�=X@ʔ߁��vB%w5�(¥q���x>�Y����K�1���j_?��:��T5P��|u�.���5��#[<aKj+���UQ�sG^G�WI����g�L�^�L���	j* ��6�/��pP��6��"V���N�5-ːr�2 g��p�m�[hE�c�vC�2�ׯ�fNz�o���v&���|���_�T{�J�L��Z��e�+ Rwj8GPi��9� i@@���CX�B�l��c�&ڂ?�f:O�C��M�I�ou ����Hd�+���&�H�!�+��bh�S'`��I�}��3���i���Md�m�4�1~S�k�Y�6�߶G�?�s1�5Z�cA�َ�,�
�*b�� (Wʤ��vv�\�ᐰ@l�z�~#ݼ�<�},��� D�黁����m��� A���W�������<6Eũ�t�)�mF�q4O������l1Q��y�#}~qd�oq��c��m)��%,�I�rZ��9$��w�u{�q3Iy�j��5x��Ӆ�m������͐�r!��]���Tã�&�p'� ����$3dW�u=h�Y�%��	w�`�R)6^Ƶ�mϪ���^���}7�s��JT�^���R���+�]\�W���[B��֕�r�À���3���jL�?$r�"\XK�9�V3i&P�3&
����<҉��*��p��JW�\+bAf�ܢ�q���D��M�|�	�1�4a�-ߓ�mĖqsrJ����`�6�
jv��̩d@�� Pa����ζ)����+�w�� 	�3Cԙ��9�N�2Z�I7T3<y>g!%�\A[p,��>�����~V��{���*/�H��ި~�t1l�1u�b�5�"����1u��
[o� ������d�R|�I��Q���W)�p7��Ŭg�b��3TN)��̤�+�Aɚ|6՘�@T�[$|�2q����i4~�	3(��71�(q[��N�p���QY�����>z	�lp-,ñ���#��vSpJ���h��b��E�ۀ��^AhTZ����_`�RWP�@=�H�2�����i
s���9�D4����hvCF�	���
��%T�����M��ҍ<oeq
�� />K�יN�>���y�l|��D�I���>�+$t�$�#oh��%��[ ��)�ً�E��O��7�Fp�Z�����<�iK����c�v��p	j:88������+��$�e�K$���G?����Q8�#S��/��Ẽ�Z3T���Ō�*q�SEX��z��⚖�0KezEV6�����)ui����Ý/>�Ag�_ڜ����^�n	���}�k��H׎��ndC�m�oB�̦��0��e�V����7�Gm� `��[�X�z|F�p�4d��rH��n�Z��W��U�3w�r!�[ʷ��/gRδ\�k�	*j����L���/LE��tF����l�l�Z߇���i$�v�0|��R��C^������� z=��J�Q_USs�Dڿ&���$��V/}:�;6��ഋ�1��2�aОȹ�˛bZ�4d,�_6�6�����
����NG�"�Nq��J�Q2F=��ݍ)�B���05��Mkfypu�ӆ���'�^���[?@#8}�x���b�«Y/f֥�PmKM��������E��	NMw����p6Mo���&��!���Pw ��G�7�K���k��	<(eӏ����pD2�&ޣ��2�w`O�B���`��V�]��+��=C@���]���p �Q�m��j?��ؒ��wU�)O"��ّ�	}���l��[��*��,��3�j䉋�a^o"s(C�01���4LD�9n/�h馞5��g�_G'��`ץ�� B�1���ڱ�}0^��_���u�,����&-��T����&IGQ���d�2�7Wf�����I�Ԫ�_��(�����2�2���7�@ݔ���H��� V%D�.��Ot���~�rb1^O8G7@�)�[%.����X�����N���C쪄�E���v8[��_A0��Q_���˞���r�U`��,���|j؀�s��F��ד�P�5��|�6�&��=ud߳�H��T��@b�|W��ځ\A�E��n� Q:�1Ч�n�[��1ؗ��f��<1=������n�'{�ms[#rc���<��0|�CU�w�&t�L��R���dW�>TDP2#Y����P��!
Jk~<�c��!�]J��A&0Ͽŵ���ʂ�į 
���^J>��Eu>zO�|���2�9M� �#y���Fn=��@�˖�� +Іy	��J��� �B,�� �e���+�����E�l���`��HPd���R4]l[eP�Y����:K�9��1���F&�=ũ���$50Ò��.Ss��T�5�/6v�g���i���� 7�����[t�~��� �Ғkf)��������J�ߨ.�#�KbF(˷�؉��Ȼ�������+<SWt%Ug�N�V	��uPr~��EY�Cb���CF*(���A������:H��J��5,��n
��X��((v�|�X�ғ���kd�4�Y�o1
�1i@���b��y�pa7�P+�[JCZ~�Iʬ�jw26���"�����o즰��]�{{ �%�o�`��y�|=9
lh�)�=�����]n�	���9�e܋~����������@N�#�k�dꇳ�g���3�H�$�2:�h�	��\��l�[���)oN>"���2M��QD����2�89NIJR�
��ߓ��T�	����UWd}�/�8���5�#�#�i�h�#���zA����k*���;P�d�9�G�͊�fiR�A�I4�p!��z��<��yۄ$��t%&�����,̧��?]H�Ě1��L��!?�SW-��$��X�^ǒ�>f�U�mW��" ��X�ā�e��LWSadF@ʻj�r��c��鼽#��#C��
�KF��k��h.:nr�rl�^CzN�C�.�E%��e�T���g���]����O}8�qc�>�^ݔOeHr��k��d�j�W�׮|���R7������zH�B*uL���9f��RLx��P�ެ�g�
�<�Fe5��aB&r���ޱ�
ڙZ���E�y����ե��Pc�J�NW�]��&K�J�u�-EwGy�C�J:�^-#2�A>�����ͳ����[�"K\�ŦWVO9ʶ��ԗ�8{�6�7�U��ĩ��23-3;m�Ý�D��
�����б�N�"�m�%lP��3�_6?|z���rL��(�a��!~j4�3O@>��,FT�e�U�f�Ǟ�͙#��7�M�!�L��k���R>�U	gE��X�0�Z5/ѿI_��0|&n�)D�������J71/�.���0g6�OWsa���"J`�/q�p\UA?Ӌ]Y*�p���O�MYܾ�n��p SG��
��|ZJ	�QN��<���~�<�7e�@�A� ��t��L����{&���j�"��F�1�1.D��b�N����?J�_��o���K��2��d/�E��	lr+�sv�+	4l�D�F�d�4��fp���0}L�ۙj�=W�:���0���y3��kQ���Z�`ʙ&twS��3n�z1�n��=˿S�V�y��S�p�D �썺	�=q�}�a�N|*�E~U\�����6�!��O���1�1����O��3 �_+�'�w��3��UC��rFE>���n��i�%p���9۟"���s4'�G �(��+fu;~	xO��^Fm�ީy �tx����tT��TE8t���T�`H��{�	\�G���#��06_!oE�:XMMr��Eh�q��� �h�vQ�H�X@۵OI�x>ȋU<�1�X_����!�$����i�ۖ.�06lX8�t��{,��V��Z�p�,2tYW5����Oˑ��x�s�;v�F�S�C3T��M�F�r����c(J��ª	��q�jh�[�9H��2�̈zT/�i�#� �.XCWK����T_Y�@k^�b4YaaGߧ��!s�2�P�(V6_�]�P�媁r��P��vj�tE�g}R��OF�٢�ܓe[F:==U�XT���c�`�&�ft4t����D��Rs���S5�C�T��i�]Y�R|�����5�����^�e� �Zս��V��E�*� ���=�~��@A`D�<�5�z��@;'cZv�m� ��\JR�@�H�;u	;=f��C���5����8=�������vߺ���|�_���#��y��x���bi� ��	le_C���Z�m�F"�u��a���9{z6�c*������� ����y)0���F(��%�xm�= F�4%?�[�Zi΀6����\o�}���\mܰ��ɭ���ĒG̴�D����C=�UsA(�����&�N�I����O�BG$�/A��,K�}&S�[3�N���TL��<�g�d꒞b�_1/��&Y��(�g��L'���dA�����t�ݥV�[�i�j����L��A@-���M?
�tU�����W���|�vܓ�W{|h~�l3=���.���,�)��@�D��e�8�8gW �6F�'������Q@'a!;�Pl��*Ţwd�u�7�.���e=��p�YZOf� �#�'��t5+&���C��N6����>�4W����dU�m[�~�ߏ����-J,���%9k$,�]�im���d�����3�i��&:@];ܣ��J�~�~�x�>~5�P ��j"�z�_Q") V�bQBD0IZ�5�6�%����2�X�c�ٱ�z��DR[�L�02������Y��2*����ϒ[x�S�b�n+.�N
)ְLG2U$6(��^�>[�P�V}���Am��[g�+[F#ӈ�n�6w��̳�,���V�!/U)-'�J��ڜ9�=�l�!?��t���I�k ��-�����0'�	j��69O���Rd�^q�%o���V;���=�f6���^�2޿k�Yۛ��!]/�NO���
��r`�&6}��1� ��dvw��O�1�W6�H�(/W�s���j�B�h/�$�k��������ɳ�'��~_���%x� ����׍���h�mp��r7q��8;�˸���ޖ�,%\�,�����U�]�IT2[�F�t�]Uc����ҧy��!-����g��IASg0�SJy�oR=����������
��?��^f��(�{�6� �A	��|=JJ�M ����9�U�{�s������U�>O��K+ ��}H�n���M6���c�����
8e�	(@E��А�!B}�J�ۦ�d�j��'bE���K�ߢ����@�}�ݰ��㤀�)���˔��Wb{���8�0��O�.��/�ܗ4vč:����ݗ��'�Ӽv��A���1�󀯰�31=\��B�s�
��\O=ϱ��߆"8���cR���e�i7�ԙ�"r�ljQӺi{(XNiJ�$��r�{����^l� ڮ�|ĳ��3�=��:�i ���П�7�x�� �[��U�N%�r�V`�V�e��.L�I��^����x5��zO?A��1�[�K����@�R�Ĵ�u����c06G�a��t��c#��� �A�N��jjd�D~j�EpP� &J��(��9���xgD=sY9���/�v ����$_f�Q���QZ�h�������$pnq֔=;'�8���1YFk23�g��D��'�yUf���W` e�4���jUY"�.'b�@qx�ҷ�Y��3�]��c���A���O:f߁|�]��S���t&�A�V�������2�8�$"�J�Y���n\zT��\r��ydy^���_ȓb��D	DI>��4��H�uN#Y5�7ꚸ�4j�;�xR5��;<c�X�w!�ϡ��"�"�Q�j��ʚ�P�D�R�FY5���L�q5n���+tP�Y
����"&�Q��c���@� x�#��m�L'���1(�}ëڧΊ.	�!|�.KR�K������$DY�}�Q����wO��*4,�,��DU���~��ᕵ��������R:{�?/��	{y"g�t4��c�3��fg��`#�>Q��8 �e�o�yB�{2sN/ S�F�������6�愕ñ*�B�S�L��'��K��N���F����[�+��4
5�9_�v+�^���\�(US�M��*�a1�V�hz����U��-o^֒�������������>��g�( m��l;(g%t�W�dye�QW
�
�o���.DT{�*VM�ɼ���a�@����J��?	��e�H��̟�J����k����Cf������������ ��a��|E+��ў�<�����C�R)Fo�$��m����d):�W̴1U�,L���t휛���I6W|�3�p}�PVRٹ1l�2�q�"N	tx62�sq�;��v���9t�_�gcg/M\>����ɧ�́�4�|GB��֨(�m�5��Uk~�&�:�0["i��ȩ8j��c��Ne�CD�%(xle��Po�|&ׇ��a�����
t��\��O�<�快���D�J���*rh=O7�7�y��n@zZʯ�[���������Z˧�k0�8$�Pwg���"%��'~j��׶�0J֖��ٺ|��l�V#6 ���1H����[W����u���T����*�5��s��ssfA�d�!�@q��(L�9A��]c�e��]�Շu���p�U�ԃę�I�Dfc]RM�I+iV>�ߧ��|tt���#39�us��'��l���ԻNC֫Oʩ���ܦ9W#�"w��)���w��@ʤ�C2���l���k:mZm�Fɑ���u�Ux�� XOrN�1����C�9�pֹ>�v;�S�=�x�Xi� ���%V�(twWw�r}��؈�8�ps���k6^s��O:V��A�I���Y(�b3��"���l��
���yls�֖W��$��(�x�j����T�%�K�288w�(���~~�7�-��Sv.�*�
H�2��"�-]-uF���|�1{�Nx�~���t���u��=ٚ�n�����@��°�6N�|ʺ��-��q>��p�����$�a!�\�(���,�$�_;�����9.	�b��dҩ��ת������-��ܴ|�{``�/_&��\}���u���h��Ӌ�3�)�W�o)]�⬩Sy�s&�]��a��Q��c�HQP�D��y�/�����R�jA�H������� H�m�]���"�ER<��xn�&P�������[I{RC$�����bc��*vU�����9,�7R�vS�#
�]L}k<�R���[��v��q��^�h�굱���� �����p�����H2���w���<c�v��A�&<��x�0Վ�U�zZ�&o��wp��2��;����+�S�ES8bu����*RL�P��*k�tD�PZ*S����oN� �~�(���^������/��J��W����s8�G�v1���p�J�?9!�X(�{�MhQ/9>c�V`P[�Ɯ��Sη� �r�~��� d}A,���Xpw&�9�E���$����S��=K!�����%�|����?��y �6�ދ��LE�~�8�w�:�5��B|
ڸ�_3R��=�i-��U�}�P�T�QWwM���}�LK"�l��F���? ��s���ue�Qy��
�R]?
yU�mG[��-U\�`���wxNÿT�`8\�(I��� t�����K���ìQ�ybr$��?��몓Ř�܎r���Gg��m���>f����1%�q�	!� ���[���O��j�H�.j�!qU��z�.�ɵ�ցv\8YŧP�ӷ��cW��d�(�H1��t��=�{I��w�42Rg�Kd�L�ʍ���N�R�q��$�ꧾ��-�Y;` T@�`<�t�f�2��+3�	A��N�}�2�������X�TE,�W�4\��S_��TEd����9nyǌ�T���|�9��EH�!���P�"�o����/ח ��wOu���8����zi�'
�u�K�]�z�<���� ���eã5ڨ��
���G2���f
�ה4���$4���\�.So�ϡ�e������5�m�j|�s�^)�5p_R=�7{M��rbÏ���@`<�ª;ӓ��iKAgw;��uz�O-��Bלa~N��JnzKYQ�r8D�Z̩��f���
ڥ#�"���uQu�:w*�GGh�o.?v�>�}�T����������y��&�?"�����.��B5�*F6��QC6O+�|خA?�� �
^�I��K�*��Q�9"�'���8���]�`�2_*9V�=�@�^�E��g����mH��RZb��(��e�F��#j�[��WJH���:�T������ʵX`[vR�,��f�e�N6eV].B�Wm��<�N�%U��wE�h��b�tf�������� =��"���Dh:�4yLpm�����9|DV���.,�mDx5;�m�t{^^t#�Y�ѽx��V�|/�`���J��˱#���KO��`@9���8Wo�@L'�FX���k<�a�(&��l9��� &' J�pRhַ��M�d�׬lν4������0�?�D���p���aW&]o�1+��	���~ji�®�e��.�A��2!�!Ɛ���r�(���/!0A-)bѪm��-��^;r24(;ؤ�c��C&b�'Fc.���)�$��H�	+fm�S�]˭z��2��#z���J:}�HH2�?�  ��	�aݤ������[%�Y#��\W��<)]���2�>D�P��Y�G���-������^8-x�A���1Q��C�ͼ��ּ$/�"z[/>��b�u-KY:��W�x�y��w����Z^$���������S�(�[bLY�c��9/��`����. mTD��o@+?Gi۫�J��Z+�>jR��x��<����}g����r��zM�ZZ"GXWe��?�Ap'X"�5s&.Yf��!�܆�+�9_�����&��58d���:&��|�L'9�� ��ִ�Z	#ߋ��鰁�����HK�M�A�_2G"
cK��ΰ$�B{��_���?�%��$^�ˌ#�Cn���>>�jJV���}�Q��!#�'%\�(�`'��?��6-D��4?��m0Ϙ��Q)piu��kg?�C��ѵ �H���	�.�sŽ�3��I�9|�{�ѵ��}9�pj��R��K��#%�-n{��Y��gұ`Z#�:�G�	�[Ӻ@q�8���\PSO��fV\<,cg{�9�^�E؈��a����.y7�*�����P�{#-��H����������P���T�6O]4V�����.G ;m���� h��0�	��26��Ì�8�$b�����D��$sV��2����hń���U�E�1h�0^i������߀�KXӌ��|�GǠ�U��X�8!M�D�����w�5��k�bn��!}��2T�]�PM�w���a?r�p1���Ή��:�����wW�<5�J��R:.)����e�cp.���V�
�~5e�sI�Z
���N;0lhVw��Y�'8¦�����O�s)#*s$
2G���l���*61{s�B��A��� �t�W�a"�%����a=��,m�.p7�)����4f���'�O�E������vS�Mϑ��4���������}��W?I
T�$$�
���G��o��uiҐ˒9ۤ��ig�u �rh�n¹� -�v3����z��s���5��*�n�W`U���@$S�����U�:��B�7D/�+F�u�C��k��� 2
/g_���0���D��]�W(�	�* �P�B�jq�iO��v%�`��_��_|r���k�O��i��)�԰�eO[�B?��4#[Lšb/�M�6�V�\P�B�PLLuى}7����	�_�?��է�F�L�ml��?a�	|Zc��R�������yck�����ʈ7B���E"x	���)�)	Ά���.���R0�G��������C;��q�%Y�R���{;�{#��jR������D�*�.�1p�C��1���Χ�#�K?���u�*t�� ��{s���z c7ؚ7VC�2l$s�B���l~E�my9L�D�I���`�5��R�fP��K<x�u���k�W|�fb��e@~"M8�s�_�n5.���rf5�p%
c�x�_Bk/;]����uv2���ت"Z^���D ���#d�-5�|�>̭3�)$��<IͭK��2��B�����V�����La�Μ���3�5�^��!�z`�Z����l�妽�������ƢXt����f����b�Pdb����ٱ�EW˄N��Cu�Z'i�a:��u��1������%p�M��5�f����q%)Bc,�������`/aj���5$��e���_rFto���Z!L��,e�<�<��/m�	c�0h�@���ť�J�3:[�����y��52^��D��(9b^���
]��PgQ[���l*�� A��ۊsO���5(��=�Pn����?l��'e��ݲ`�X:˽����$"��0��vM�f����:�Q�RŦa߅�i'ě�1u��Q����H㗗tQLm�IY!��<r ����G͵)}?�:<Z;�}��~����91�k�'�@c&[�w�X�c�z�Rk�0��,b�[���@E�8Yq�l����(8<f<.���)z����}
��--��H���$HM"��L��n{l6�/��?,�"����� W��� �}���"� m/�n� ���.����TR~��y:��O�#���˷a�k=6ޯ����rV速���H2s^�0�:����FO �DR�.�/�:�<rY�i��w�zb���x(���õ��5G�s�K�d*w��:_x4����%��mK�O���@����V�n��0;v�-(�2�N���|$b��v�b������Ѡ�-(�Ш	���9�!BfSʁW�Z��7V�:S��^X!gi;������x?M
�?�ewJ������@�����=��ΰ�#?F�߱t�y5������cq����ʤ]�R���wTY?a�|ۡh�u�_l�V�K�r�1rzQ˂��A(��� �$�-�i��(�8os݈i�31��4�����(qt����RڞԫJ��<�Ɵ�`8JlțԴ�x�xըh��x!��ڿ��TC*�H�?�d�$dU#��WLO;Fr-�0@vb���'����:�����(��D�����x�M�O_m��VI>b�fB�k($�A�yXs�� ��l�T�hSWQ��b�V�k����-]���<���� �v�X'�Z���%��*�,�6�ۣN>m��XcE���u���)�峳.�E�l�x��Ik�޵�l�!�l�FN[��� ��+����N^��e���$t�̲I�O�z�m�dҟ2p���
�ԭ�JF�oKp�
�!��0�S���}�w-�댉�5�"�By߉�ӟ<�I���p�_~A�Ճǰl���HE�/4�rS{����s�6��i�ڳ����ɏ�~a�p)�(O�ì�=WJ��W�ڸ��}�U��+�A_;K����2��]b��ɰ`�kt��1	�;��������̓L�_��<�-��|9�:GPf�͛BB��G��H�6/��ٜ#�<��d�l�T�@��8ez�,�`%T��� �K�
U�4Ӣ!��ajl�7�K}ڋ�~#?A��L�4#C!3Z6���?v������)����e��А�����x�����`���p�����W$%g�\c?t�����< vN����zXC��810ZU�v�����G�����l�/x��A��jv'&�oDWO��P�`�3i%�I�f:- �7v$����rgh��W�O�/�h�|�V1��MZ�a���|����֖�7�L��X��{�^�� �v۸�8�"��?B�L.O�]�Ȯ�E�aD�{F/ZB�Z9H�'NF=�t�m��/W�M����tH��n�A�Kg�>���e]�m���7]��?%�GB�2M��ó� β��*:7����+��8��w	����}M��|�h���5s>��_:�p�5�c��j�>�B��A]QX�S+
��X�յi6X]�M|é��c���-��+���v�}�Z�DN.N��> �Mi֖	V0^�޺�D�:��]�����w�#��(";�2�x�[��xh\͓IWּ�tiq�ё��d����hj�i�4�T�Bw$�����WZf�@���{�D6��-Ȧ�=8� Ĥ��8��a6pm9B�A̾f"꺤���+/"-�qfQ�|ى���6�+��7y0ͣ��	����yO��[ $�Q���o,���.	�'�{ٵ�ypr�_���,���0К)����.���5$v��*�!>ʾ2��9-�X��R�@z�����]X%��i�@J��0Uu4�[̝g������Zz�@#g�SsC�.&��}���.�����^��o�[�8O�-L�!8_^X6*�Bz7� �K��r���CA�a,gĽF���xq��m�kQ<���O5�'�jSGcO8�^�9��DҺ8C����*,�ɣ"%�&J~۾d���=�7�c�yBnl�Qe2HT��ѻ~��Y���>7`n����g��l(���-
_Ps��b*�&뀗�+��9]:sT��\zK��U��h�
��)���%�0T:�`�?�c~�GQ���u�{@�lco��ڻ�����p���K�M��@
0]%��ϚW��72�Hks����*:V���~AI�*��[I����9r �HD�}��`	|1��6���W��߻ĩ��$�F#N��ݭ�{֢���2/��թ�'�=�(m�N�ƪrM��&����P$wٟ�}Y�+|���Ά}���;�wUg�a��Y��<V���>�*�k�V�exq!e�ÚC��P���n���}�O�{�kj\�S��R�.�IR���c*>dqI�-&9<���*�`ć�@t���ݤ����݁���Eb�ȷ��gU�����ʤ�(e�]�F�4y��<�|m����'[�Qa�Xn���(�h��HOKͭm)�O������m!��9#k�������c���z��#�u}ɓ�\��Cz-u;  �w:V�E��f��Y@\l��M�k�'���ur�a��!9�r
�d+�7���f6ň��|��|g$�h���ҿ>&#57��]|i��d}������ϓ�8���#�w���+f��/�9U5��V��ӓ����*��}�9���������l"T�J��Tbn?.��j8�PX����6̲Z8�tDk�Prޱf����~���\�%�Qk��V�E-�͂;c
V�n����ҕ�m>+�t�e qq�B'��6Վ���3�˶��Յ�z.�����[H���A%�b��mQ�t�l�g�[��Sx^��6E(}*T�>5|�ܴ��&�:	�y�״���
�鼺�T�dn�<�&U�Y�Q'�ë��d�5E�Y�x�M�p�����V�7L�C�ơig�u-�i�.Ώ���\��Gu��b��58')���H��+*"�~2�,���veM+A����n����->ҽ����u��}�HI��H�����q�q�3{��o�<���{������=o�m;�s&L��ݠg���b���𶙅d��:I�a����pDҳ�O�u�|MPI�El�i:R]��퐠�e����;l����tHi��M,;��g�Ȓ���j��No�:ЅbyxlU����6�ѡ|�d�H�7ϯ�m��$�6�{R�I�&d��������?P�B���	*����IZ_mP�i���g`T*��%��{��?��M���P�k+�b��ծ[��j��sRA�B���%�_�I�@�E��\�C�K�;^�vF#�E��#d-�xٹ��kR&+����?d��<�Ŭ5� �=f��:��IgUU�m�Y�����`	��!��f��DXg^������NKn���͞�Y�@���DC��0%?v&r,�Aq�.O�\�Y�|m���� ���|���h���{��b���\��x�v���Z��I�� e�T��t)jB�������W& #&�+b���9ws��/��;�R�����φ����p�^���yLru��D��r
�k�5�\�}����]Oji�Q,Z ��OY��ন�ջ�>��>���Tt�N�Ά��/�Ѽ�J�?�Y�&w8<��r�g>�'�.6��f�q�:o�i���A��0�}8o�Z)eg��o	׮�y+@~q����X��[C�����	�&�͐h�����(?��E�^| �KY�X;?�XN�����b)�����N]8�+P7&�.��.�X�5���W�e?�'|�}��ݏA��7з{�_�:�>���}���(&G�B�(���V�d���>���.N�q��6n�^|�.�pn���c�����ފ�l_ �sjTþ<_n�P��r�o����$O��TLO�S�"��G�	�~3/{p�sP�(�
��l2�h@��*Gi6�NW)�?y=�F�p�}�m�E����#�0=:��tT���#�{-���L��r.۱����6E?��rdZ�sMP�b���x�i�X�P�U� a߉HA��t���m�pG��KŨ1_�s	�P�{��8�R7IV�!	5�t-�@xaq!p�Ti���+Z��yy�t�j��*�AGܘ�\ۭk�Gi>�W��P�4��X����qY�7w��k勞^�<�>��>-�t��X|�!@����]�$=�kt��W�߸fئN�-.A쫄N���le��C���^��ݵ~�n��ʸFl}&8>,�5�t�0����;�QJ�.�d������+�%�`2'R����׊�Ḝ�S�tw
��d��S�M�k&���d"2	�M�~4H����k�ǔU�i�ed2K����s��bB�EJ������	�S�����<@��tZ�ȴU�U��?<�M�|��x�~�Q�ߤru��9�~yF��:p]{�y�l�3�+o����x�v8�C�A	�0�0�uWa~ �61�o˃�E��[e�opy�dH��^��ݶ� �$�,ǔ>�d����5t�9���ui�x�?"�G��t���t���W��Jw^,]LE9Ք����ّ�ﷺ�[������
�`s�%�E�0�c�=����̑t7@�^~���$���]�r�?�i�����}�� |��O�Tq
#���Ѭ�5
r��f�{2�Y�@�؟�j��⪄���w�Y���*�Ⱦ�?�����v}������8����Z�+"�7\Aq����+3��V�2ܭ�-.�e�q2���*[��B�x~"e0�� ><S)�$��Ep���}rA�/w�1�ViW�)�ɹ�D�������rr���(�?���!K���&Qz`���*�¸&'��G���w��A�Ss\i�^�m��.8m��a\c��ʊk�d��>��������[.�c�p�d�iU"Y�%G�6M@fU����M�l6��d7�w�l�?�Q�M�ݨ����x�P����t��CW�%��Y#�D?�k�ҹ%Z难�{�%�>X\�;|a�]�.<�#Ph8<_ �����W�D�hfO9�!�� �JNo;��[}W"����lpIb�,��\en�B�������c%�o���Be����s�I �����bʝ�;e���cc��R�T�5��GeJ#��F^��ѻ�
k	9c�~j��dA}&��VsD��=����ڨ..�n�w\(\�G�
FB���1
�[#�ӴB��~v�t����zIb?�F�3,B�q�d>�T�c&^UyC�P�>�h%��o;��r01h!`�T��M:���0��w[�
 <�u��0��J�R�=�t��F�Ĥ���e<C�U�(�-��W1����*Q�`F6
@T��C�0N	�Sm�\�����i��;&�����	��Z~M���@�]$T�a�^��PE�%*}�V2���ͥ�ݸ�,�\���T�,���?M�-��򜽨8��J��-Re޲�Ɋ��6�/�_��D��Q�ڢ�M��/�HV�{���G���\5�]����q����za�S9�3N�Q�*���}_��[���k��r	�7���S���X��H���gU�-|iW#PO�9fO��<%�X?ES��y��z�&��Tm�7kZRt�_�����ƕ|��`�������Z���I\ʎu�I�!R�kv�мZE]C	��6�P��	K]_�����������l�@���"��h�H�C�j4H�@�]��?1Y�U�O�Wr�u-W��ݵ��4�yRoj��4[��~�Xȯo&����Z��\�}:j�� r��6 ��:\o���͖�F��b�1F$�P̒��8�^�����䰇�
U8}�URt���G"4�~�1����֢�M�0��[,4�M����o��8X����]��{��d�J�Z&����7RٺF�f�T�9���ɨ0C3q�å��t�w�O�����Q�CT�ĉ�=�@���S+��Y�<
��h�Ł�m����f�O�4f Ě.�iUI�� �5k�y�%�O�J���IE���v�J#σ�E!B�}��^4���n!nP?��k;�UxM~�nΤ���Df�&^`��V��[X�=��@���_=��J��&���'��"��9.H
����z���Ώ^V�Fi ���Kzo$���u��N8�����%�Tˌ$E�2H�����m@"�_�d������Ő�es�(�~KE.|��d��E=_�?'H�|��o����3��	ߦ� \��r�7;��g��G�ly���	�E�le���뺐��D�*��а�ij�4ha��P�[������5����i%�Ǜjl�O�;ͦ�U�3��P+ˑ��X�|���&Qn[	N�2����[�H�a��nAցM���^!�A+�^��� �nqa����7�X�6>#u�;#��/z�T�{������#!��jkItP��.p��\0ƶ���~qo"��4ޮ��ƣAV�+��!c��o����d� �J�D��g��u8��Nu[�Sp�yy��5`;������ypT��4d,FH(KP�2d���"?��ji�Ϭ������E�Y�����a�<�k���[{ֺY�ѻD�X�h�K3��� �,��}��������âh�&lv����� �d6hC������i��_�7�`$��B:��Y�;���g��{[�&?ʖ���3)�Z����!&�K�/�T�'��e�?�����&9�
C/� a���.��&UL��&6A�J�s���]>���G��6��,�ꈚ���sKc� 3�E�lf@��ˈ��#���3��ߟ�0V��a�$��2:��S7� 1�m?=~�[�
�<��|\��:#��v�! �`?1�A3
V�`��W�l�<b���T0���Kʞ,��f�}����7%UI
�tq\�����ja�`߻�~C�h��MT��O�Ӡ��O�C��.Y�t�u?���u�d�XՏ�����0	�B�(��6Ų5fbʓ`yc����"�2��԰, ^uH:F:��ᢚ5nV���@��8����y^8���V�*�\�TT��l>�=cK��so�G����B�8���D4M�Gŗ&���_�S9���U�D<%OJ2�
������-�1��5{`���J�u� q쇁��7�_{}a�و���:�L��Ph����o��4�+[�n�#g�U���C6Zq��&�:�+�-^o�A}���2���w��D�G8"`�Pf��I7י���fn#`,���F�z��?�5����<�4]������l�1WL
7
G�Ā}����#���0��	p���s?���!�Ԃp�Ǌ�P�P	=]���]YQ���/O��(� ��ƴ��f- g/�/Y�����e\�䨨����Ċ0<؀���iD�w`�dla�(���׭��P�7V�fW��k)A����0	����VR#цp�*�a�L��4��K�0o�ύ��/��kݚ |t_�
��(��K�6�ņ�J74����{��X�wxO�t�t�B�%�g����h��4���J�&%�ߥ�ǝ&�+w�ъ��d�fRQ�!\�L4�8l0ii���;Y�q���+�ɚj{\�=����!�w�waT��><Ig�BE��C�7R���9�|U�9���䚑�2R��/+ 3є3���b��t
��(��xiq�{J ����>�'ew���n��A"f떧��y�����Et��_�Z���>n�Jd`L�q�K�A�L�x�;��s�E5&J?,��w����`��>�a����{�Z,�LV�8}�������H���w)T��l��}X'��]��QO)Y'_0L%��0��TX��S�Wcp�����e�	�|�,D���'S�v|�ՙ�:�g$��@X���)%��Mt��Fa����w�|"_<���o"?��"J���Lk����iH���J��`��O%�
�����Ƀ?�9!��:���fmv���=���2&���l�ky_��}��C$�m�8��?uq�d)("?Oly�ԏ3m����!'��y=�}�3G�����t�L���O�؀=�.�����Rx��Ί'j�� GI�O����ۉ�o��.O�Ӧ�O�k�C���e�p��أ��f�}`Z��� ��X+�(�ǽ�C_�-��LIZA7���xu�1R|���j�*�v��@���o-�0�{[�xԃ{��e�-��1�d�������46ù�v�t0*����ӷ����������e�e��c$��ͣR�,�C����G�4Za������t.�������D��I�<�I}����i&By$N��}�~:k�M�ݗ�#m�v��la�G8s�֫����c`�^��Rݮ,Ӝ')6x��^���z�/<lyR���_�ԋ4؄6�Giu�+�/EL67�f�&��_��:X-��y~�K��� M�t������P���j�D^h٧�
3̢`$I��w�g�D�.�+PsR(l�;��������oMD�羊��"��EB���q�Xy���<��Ra�e�F�ޣ/m�s�N��a^Q�<��o=��a��.�������aպ�8t�%,���w���� o�R��ز�9�p0e"��b�Q����r�4�/6��P�d\+�pYnU���>�J}`�-���3Ǫ��C�tJ�>�Ay�~����L��c�ϵu4�����Ǭ6���l�����t[P�2L��+5��J~��΍�S+�ݷ�3�!k��"�8�4�L��-�,D�v��drdM ��~����ً��$�4<�����:D
���$.(/�E}����^�����J�ݼr�{O�Ξ��^����r��=V����s�	+���ɹ]d���9D
�-�7x�6a�<yAr�)6]�TOJm�jU�;[�]�#��L��^��� e E�H��Lv�mJ�)�Q�kF��D��tWLٱoŦ�(�RJp^`�O�4&��ߠy��`ճ~C�δ�N���pF�I�3�\Q�؂yT	8�|�ŋz�;�"ph��BEu�=���<Ys��f�q��y��J�����.��RB������鲶`@X��ڮ!	�XY���3�*�r�\�j\���:��F��ϸ_4i� @u�Y~o��-"�Z7
�Ic�>#���m����K��%'`T���1N0�vUp��Tu��4�𨉝Wl=?΢S2�,euv�����ʀ�74�fw�d�M�B��??����	��ε������9Py�|Hq���S���Z؛fTҒ@:�Ԋ|�m��&�
^� �=�P�iǱ��sz*��@��GLN|th��x�QƮKݠR��%z��9�����2���a[��* �L.�_b]��Y7B�_�X�diy�<|��S�՟ܨrK}h�qj$��v=��E�b!SR>~�@S�B$�À��(S��H��2p�a%�uʧP*3q��:�W)z��<*n����C��;���8t������Kw�A���-G����6)�_>#�����= AٺY�`����V&����Շ�֨���~�!��~�Խ��Å����D�H��ч��h����I�5�޹��Z��{�F��]?G�l��F�������2��~R�}���/�H��4�Ƥ�}7��x� ���|z�"ӺR��TK;���<�����Se��s�S1�\�!��*UyT���0��0�O�=K�/�喉��m��l��ɮ�����a�䟥7c�S@R�u�b�u<g��� M���tU@#�>�n.�g��˟UN�Y���w�F¼�70OZ(��Yi�]NjBV�E=[����W��-�v�-B��p��҃�cL��,�z�g�b	?c���j�����N�ͪ��(�KA�^3�ȓ4�a�T���H��")�<����ٲ0!�Ae�i����C��s ��ۓC�"Z1 r��4��$w�i���t����p�M*�6ZߝS��b�z�L��d�IZx��� ��%%J}��I\
	M��Y�K��� �q���9�$�Nkn[_L�X�w@P1mY� 7�� �¢��������f�`u��1DJ�k��d��Z����|1�ߋ&i��C��&�aʅ��������`'���|Z7����~�`�N ��=W�⩛Y�q�:i�p��'���0N���#Q]��qO/��3�8��?c���\�����H�%����\_@U�@�~iH�3\�Z4+#���.�pUB��A7���H�"��;�W�PޯKC����ʠUY[36᥈��F�2���.�7�qI�Qc����8
���E�h�9嗬;��ml$�/�}}�F���V�H��z[h�O�\�ˎ�3V��g}��ȀLb��|7��8
3�U��S��|V2�e=�:$*��0�����NR���^�ܔ����U��i��B{�X_�Z2i�[�A�p��:��o�h	����SD�����l:;?W�^�y��I!���]�+�Z�_F;w �Y=l�nǶ��
�R���b�1�=1���1q3��	�� �T>��t��*�2����P\��;@��Z�"Z�4u{q�.��}1�bH�W�o"��E�(t-���3���?#���E�l𣰳}��m��o� 銆�{�h�7:.���4Ql�C�^ �=��a�6f�DU��̑�-��z������ҭڛS�C��Z�k�P��i��R���g����Y��f4U ��m���2h~A�܄�)�hT&���,w��:�D"��P���깹E��c�B7��t�\Z��B����U�S���K^֑�[�v�{�X\XFO�?�,���T��=�V��R4��͂
�P�_�hm,ط�*��&)A�v誒���@K���˸j�l5A��k��ބ��(��Q�!/�TN�lr9V���{��7K��i����wѓ���k�I�sZ���A�C�aPR+��ZI?�)��n~�jp�l_�V��;
�c�n'�2��(�&(8�X�`=�>���(��i�����o7,����%�͔h ���C��>`S-Wm��Rק҅�qo��3}j�{���N�&%��s�����WL�A�����)/	i��zd;�&@�]"Z
0:�u���~BMh��OŻZ�B�]��r�?j������׋7vt�->~IH�
l��op>���*��0#qBs��G�,����[!q��
�\+�\��r�4�"�"=����e��U��;$j�[�PlR���1�	��^���+�,u=�LR��C:i�Mؒ�~-��0��䮬op �H��[�_�)A9$��أf�s"�R�s�F�  P=��FHLl��Bh(���ob|�_��~��uQ�8��
��Q�CpEA�~���%W׼0�m�6�.P+9�����������G/�|�g���ʚ�W��IxV�A�l�c��RX�,��1"�\�E	R��47���]}2?�=L�ޢ�S�A@�����
)F��>r��ى�ň�j/�re��;�r�����3�:ݡ�� Ą)u���ȱ!�5�F[;P�����h�A�>"*���I�A���=�?� ����Ӱ�;b�oau����Ó�<I)��6Re�4 Qx��jd�x۞/��1F��M�˾C"���0�51����H��s�� 4�%�Dc��'�m#Χ���C7��('��U7����h�Z؏@�V�	K*�3e�<M�O���S�_�t�'�����R֧ x��QJ�� ����g~����n/{xP�~X
�Nd��s�-�s.�_�]S�5(� ����=�L�9�bM��|�և���8�?mH�ݼ';�'�B� *"\�(��gE�Ƴ�9%�`4��V�M�ښ�+!�(Ho�,̍({IVJ����K4ŷ���w�/M�=�ߘ[�L?zu�̷�1�˙��7���P�q�C��V7�A�Cgva�O8{eW��)$�� 4�:��;� �����i����Y�b����p�<��HLJ'b:��t0�Í��iah^�evJ��c���1;��ਅ~D����"7�`V�^�̠_���"����~�F�;1�h&I������^�B�p*>��~���d�D3�s�7l���F.h�����ό1��A����I�2m�dAG�c��in�S��jʽ�y���ca�l	���e� �P�5M̘ϞٛP�`���j;T�5u�`,����q����2��
��B#�o0l	,{M��܈"8�~/ ��S�2��Z[�}6U_���(��/�]������%a����P�ʎ��/��1ɟ�?���Ob2;�-dٳ.x	��=;\�ƃOF�g�zC�1̔$w1����l�����B6�}���2ɢ���96ǵz�H���^j�A{� �X�hWD� �,v"��ohTA��P�O���=���Z���v���˧��=�$�W1֪F�rǺE\�8�u�tP��F�O���.�}��Sh�����b�W`�ZC8k�ma~�"��Ȯ�!�)��uy��,~�ZS2|�� `G���gp��Ql�*��˪��ܫՏ�������5�(#�%�= �Y���62���.��*�ئC&�ӯ���4���I����!�k���z����l��}9�zM�ٿ�$���~EʓVa8�_uI8}�Uo��/�]P��T����=?P���?�.�8���΁�a����*\�Mȋ&wv���n
A~�fx]��άg~ಳg-����"׎�Һ�g��P��<鄸�G�?�2%K����B7���b�+��
�����īC�A��;t|^s���=R�.�XmE+=�?�9�A��TZhð�Nѧ���a�:��"��8&�j^�Z�ŧ�%(99��j�K�Q�^i���#� T%�ơ s����&Y�09!l&�Qk��@�D���x\&.Z5�7z�aid..Bq������������Y�gB]�۵���9�PQ���F�U�v�C�ҁ'�8�G�e�k�_(4�r�����9���]I�_eI�_-�K��(޾���WdE�~J��GT~�d�����g��tLG��2N�{]�u�����vV$׽����i^�ʓ$�ͽF?f�������H���Ӏ|�E4x�����2"�h'�h�j���sM�c2�>^Ih|w�C=|�f8gh�v0�m�`r���	ۚ�>XB	�i���-�X���u�V��q��(*��`�V�����̪�C����-_ ��d/c�\AK^ʫ�^ �Op�j���rgB�+ʛ`�e@j�����f5p�]d3|=d���u6�Q����'���X���r]�?7� �N�j���o{�:�4O0�}��� (ƱAKx��?��z��VE{R2��~_�G,� �	问����?ɶ�nh���d�34�N\����JD𢸼wV�����"Ϟ�����g>�ً(B��ol��[�kcC/�l@�~���p�tu�`"t��VJ�jDj1��8~��1�Ռ�j*�<411����lC$�I={1@���	�<�b��A	��/�/&��G�cG�ebo�ȯ�g������Z���<�M��&�'���>t�!c4o��GJ�Zgǣ�h���  �L�g�V���\�DlCI�D���#�Y�q/�I��@ޓ\i���F�� ����^��'t��Ii[ə����>�N�*~�u�N�g5�k��EHApV�t�T�I7I^���'pK�%��y��$#��!��x2���.�}}�U �
�W��m]�56'#���� ��[D�*Ĺ�z��щr��c�%R5f��uo������C�� *��d�m���J̦��6�*����d=���t�l�B�'S�K>��l�YBׯ~���a@n}
����ݾ�Ԙ�3|���0��@=�����\KV�/�l`��Lu:��J��a���}�8 T:�: 2�i!	i�AҰ���u��h�C�-pl���l�G��y�d�|��b��j`B����V"�5�k� S6�4z�'��Š�_������8���9Jb:��섊c9��Y_ �a��Y+��CQ������J�ha�<aNe�Y}^P~[��.�^<�)�|�s���Sm�N��,���]��D���GC�p��X_?�_e�w�kJ���)p��f����|c>���C|L-�@<gU��{���jfwK��:�"v�(%�L�W�y��^� :l�,_�fW�g��~�-�q^S��y�\�Z����]�9ؾ�J�:�Z�_��3L>��iL�d1�%�6��$|3�j��8
�bh9x\l\�ˌ���k80����]���A��`%CY�eB��7��2��o�����Uē��۳�8T��:�+�.����oVM�PQ)B�=�4NJ�xһW �1�D�%���FQ�Fs.��|���z,��킦�zv��X�$���K��s����2��M�W��묃3��KAaWk��x�a� �}s�O�ļ#ܝ�7K������%�F�ؤpnc�_�SiS�-�uun�:Qx���Ǟ�9��Z�mW���]s��֍/U?��BF��}���h��<8���5�� �H��<�d|!��ˍKry��&�3Zc��ԝ�(���8��(�I��1�F��1a%���F�hz�쟨Cr�W%ȍ��X�/t���RS���ag��:]�g�Q���(�h�`��x��F`�����0�6N����U��L��*�;�<~��ȡ��K��R�W�糾�`�g��q�\�?��F���J��*E�G���z���C��Y��E	���O o�ss}����vϋ�	�(.��Y��Pcr�PMK+�&�):��	6\��L#��}K�((Jc��]5�^L��1x4X�vU
��_A��3`&[S�V���-�H���i��wC j���ZI&�?�&R�7�����pN��a�(qc��&\�+��Pb���=R4�O���m��9��,u!���IۼB�R[,7D��h�H�����k]��J�l�u2�èyA�ܭ��wF0C޸ǽ��f����ɴ{��7�C������[^�8����؆�6��e)Uo��
���0�u|Sa���y4D�̵�;&@��}?���2����/�B�lËC���d�Zb�Po؝����O4����#^O�a��
���(�WŢC!.R�
Zv�W�s����P�;ҧ��9�me}�h��t:}?�nxf4��<�2.79��/2Z��ӡ��Zk�	'r<a_�̓w��Ž>	q�}2���7\鋒��������K<�T��J\ͭ���u�q� Mi����P�٬D�֞83k��A��"^�� l��n�64?�H��{aegH��7"ev�|Iޢoz~��y	KU�Y�j��k���6���v�ݒ��Ee�)�i�w
�M�U��P_֕�g�`i�q?�t,���$0��>�xM`�	Ϻ�i�5��f�%�Ϟ2Z�9Qk�.D�u�u<Q�d�ۚ��̹�[0�t|�÷d-%��|�h�����"��+tQ>�إ���ւ��4˓�]���k�G�8������IG5��l��@���&^ 㪁���em��be1E���@�����w��Y����b�+�j�.����Trn�F�ˬ��[ж�}��.���{��]4�!��b�عr�G�^�tt���8C���C�����;�Vڒ�՘9˘�"��>��v�.�k|ߙYy&$���̩�X�K<��aa.����(�?Mh�}�N.<@^������`�$O!W�`Cb�*�Ed�و��B��c��37�,�!8r>���"^�uV��6�(�����T�� C'yA[ts�����]+�s`�e�wX�<N��J
�s+�S��*G���|��g~�[����T��ui�۰��P�ґa.p������7�@�JYU�&��U�)r�A򵬒��m��F˼�����r=�J ���a�i����c;ס^���Gf\QO[9�(/P/�m�/�g�BՊ#G��W�6Ƚت(�K��)8؅h
g@��&lq�����C�1�����Q~{�凴!��立h�j
�Ocy{R��~E�+�-"��ۑ����׎jy�xDب,�)<�/����{�̆=�2
Xew�=E}(KO��|;}��A4�<��1
���ة_�ڠ7F=P��S����j1	�����P:��-Ym�f#<)BV�I�a0�{���{��!���eh��Yo�yM�F8�j��'������ת�3�8Xkv��WO���@Y.|)fy�+K@x1A�������s������D�5�+O���e-6�)b!�e6D�I�5�������4�les0Y����� �E������g��D�i
~��bq��V��/�)��g7�O�N�t���$k��l�/��ઐ�LŃ4��!M����̖М�E���ٖ��$��t��B��K�0bQq���tw�PQh�	�!�E׊Wr����d�� 4�qc�v�ҡ
/g���F^Ƥ<B��X�%@M��A��?�I�[����rf+�%��#��F�NI����yU����Qd��<�����jDG8�n���0j��A�V5������K�U�
b��8-��Am����)���_�u�n	F��<�d�x��C�,��6�^A����bݺ�P�D��{�;A������#H�Dw�~{uF(����*����/I�N��o�#��P��Du�����n�֘ ��Qظ$���X���$T��͸�5���\�p���ɒ����Q�#� ;"�d˄��J�mi��P1�%�������4S+@)K���y�Ѯ��C�][#7p.��ꟊ��� �Opm��Ib�H��n�Xm+�"*����DŁ�w�����`��T$L��n᫛:"BG�r�'-���q�=����D�JLx�bďhI��s.��嶇�5�_J�����f\x��Φ��Hg��8�g�$���JPM���\������"�3L�p�X�]urw	?���{#������B!0�%�4o������^�)��SN�>��%�8��L��#�X�k]�e��C*�m��G�Q��e/�:���E�����˘�F�c��-G #�]���ࡾ��0��:������
z
�۶���_��N�W�j������l�.ce�UEi>�Rle搦
��D9�����Iz�(k=��q)�y�4j(X�Y#6eL@��T�2 �Jx2�ޠW�����(	�y�P�� eiת+�y�b�}����ͪ���
��u)�ؘX.�(>����7m���{e�RtE���ϣS#�<4��ys�(z�\l���X��m��Y&��U|�b�r���h�'����Q�c���c����N���z�\�>~��F��)����������B˹��RtD��c�7o�<��F�Tf�|��-oi��b���b�r�zZ��G�H�a#�Eo$�X�qWac%�]6 ����Z��ެs���
f%a�i%G����&�{��D�̓~^p�Sg����ҡ�8ٍ��ћ������;�� Y�.T4�.�YEZ5���h����r���?���1�n��_��+��� A_[�'.�\�Ntl�ј�6�ed�}aR���Z_S��"V��(Y�Jy��^,����ܙ��8H��D	�`�2^8%��/��_���(���onm�v��dA��5*�4�'Lc��N9*��`���aB��i�Q]$��7��x��+y�qj�i�0n���H�<f2������LЏ�U?��}�l�H��������.��\[3����7eV���xZ���.��(�����.r+s�S<	��|M��ﾸ�&P���w��mz����i�XMU\���&�	#(�^��e$N� ܾ��B��T,L��*�WZ�.ͱ�XL��e�#u?_9=n�_c�Uǔ��\ڸ�������2��v�<8����Ƈa/	�Iؤ˽[��	��$�u��9Z?'�/�3�hZ�8���C��7���~}-��@o�F�t�-	(jsޜ%���Z��� ����[z~��re�����
��j[�V�ٰ�=r���]_^��'Z|s:n��ua��2��"�@ �W�{����_�0�4S�'�u1=ʕ�"�5�xJ�m���eJV5ea:�����w�����"�W-0d� ���c?�C�*(��B�������*�;��p,%�F��2��UT G�D<Wl�.��A���G���Bߜ׶�P�o�04�93�_�0�ۜ����^�^����i�3��`=�s����`����HI+S�?GG%���ߌ0t��92P���o�FЏ�k�-RG��2#�}�J��KՉ]$-���������@��#��rI.V3�r"�"C2�.F�F�%(�[��@:��0���C�ġ0�E�����_��,-:�2��v!�C�[T
k�9׎[ң����U��\��E�\�~�-�h1R׾R�{
Q��R�f��MIH��&�?Vs�MG��������;�zj����R�S+Y'���$��3��_p!*���C����@@�j��1�(8H�d0��7(�"ψ��x1�i�L����ɟ��6� !��j{�JF��;�;D����;%~/�5�3���~�US�G���Rڽ)�KaZN�a}˰t���liK�B
XQ@WH5�:�"קB\��b<�|���w���\z�i�b�=/��\����}O;�Ka���C�D5@��]�xp#���O^7_��b�\���}�o(q�h.����ȗ�VɄ/��.�����!�����V�o�|j��1c�N��/���:�X�)�(\�pÁ/���^mnш����f)*IZ�T����8zP��8���|t*rC���Дe����ŭ�I~["WI��<4(�I��8��nK5Fx%����Օ�z,�O-21�̋xN]��{D�-N�Θo��u9m���7lE�"���m��HW+�o����w�����l�A�
-���h��Қ	���jFMt,�`h�}��:t ��JC<7)�b~Ro�z�s��γ������Z����
����4���&��M��]
����A++�Hf>sd.��B��ʙ�=�E�O�ĝr�ψ��A�&�֯{��&��ąф�p-D&ϝ�d����VQ?�����^l#��s���'�w|bG S���n���g��o2⫿� CL�à��z_�pQ͛8y����+w���Iؿb���s��ߑ6�+��U���KQd����Zz(Df��j%e����]V~f'4'�O���tĀ�u�x���c���9�]�H���y�R|�B�#)�)=^�AH���}G%a]3D'K�#�J�ܧwC�\��Щi�ԝm�C��5�r�/�z1��V�H�6'���.?���m҆���q��`_�;#���\�c��bؐmVr(��sS]�O��S7P�e�����Dv��r�$�� �@��S�蠿#�+��|�� �dƂ�Sn�>Ot�i�%Y��*���9�-���.Jx�d�U��e"OC�TpC��V7� �l�P�*�����Mü
��$ ��Xn�x����A!��̟�P��/%���d��새�D��V>T���#ȴ�1D~(@>uɀ�z[Ѣ�q��c�-���᱒�:}	�1�մ�MK:�E�u��'T*]|dv#|I��c�u�)��`�w���i���0�zi��+����7`r*fO�I2.��.۩�B�Ɠ5���Џ!�M��)�A���mU��^ %�x���t���J��-�4ϱ� J3X��_��́<4��a�����piyH�y&��� �m�~B���"���B叜>�R�yg�$����.w���kC�l�D�8��4r��X��ь�υ7"ڈV��#A��h1=	�4n%3�mj������c��ĻB,���s�Xy�6MɡZ�_�~�ͩ�+�w'g!�OZ���S+��
�� *�?�ݨ���1��̵����ŝ���v�Q�G�VyZ����ä6�,�{]�����oG�U}���`���e>���Y��\�TQ:�Z�H������8V��skӍ�8P9VxV�G|�m���/X�i���Q ��=�n~�Od�3��b+E�K��|`�iӼ�;�@�����w<���H��9��:%��g0,��J�Z���瑆<a	�L1�UyI��G��Kg�!�2-'��b!:%�s�m@�1�빨��eT�by��F���ތI�&6u��]�=oPs]�^u�ZA9ܜ��z����d�ժ�f�#��~��IkB�::�>���,M5��l�&���I�"�o��7�ч�F�&?3�!���c�4�h��E��C�
���T�ן-�W�����};���q�x�poh�-g�X:BbN�z�#�d���1�s��X����ߙצ�
�t�а���D���\WAf�x�� c6�ct�ܴ��fL'*#௼e��d�)f�J���0��o�&c�o�<���|�'XL����=b������wg���H7���v�jW�'h��H������{;6���|,@\�4�pp^|��\	JL�XӒ��0l2�)r�{>��q;�5���T`��_a��9�ެ�1���t=����X7ڌ��_�G���X�o��J�j�a�O�gw���{��_�0�N]�?�"*=�2U�)ޛ|=���:�fQ���0�x�@~���N�?�KЏ?�右�bh�@��F��s'b��;J�9,[ۈ�F�'��C���^�Ѥ�\���ڷ~�x�+�)]Bd��:m㮟�k$�!���Dj�ߐI�[��θ����+��g�p�����Ĵ�
?_e�b
DC�-	�?G��>cP��!+��]Y^ �g��:�:��p+�w��>�Ya�[�ҽ��1u봇*5$7sQ�{y���t~�5�d��`�%#���gt]�LY�R���x�>�@����4 H(���
J����L)D��k ��W������2t-˦�W��j{s]2��Q�Om���������~���to���X���]`�l�C`=���rޑ�:(I���P��@b�
_�uH��a�_ ��n�9�*�	a^ ���{ϼ*��nZ���9H���z@�An����B�M�3�ヒ~d�%N��J�s�N�n.��MHp:������2i�^�NP�+D���S��a5�'K�Z���:��;�J�{��H���\I�X[L	�5`]�',/X�@���R�{v����Xd�[�T/9g���z	�5Pϋ-o��E0Z`�}���E�?P���B��!,0�w+����C5:h1%��^�e��ݎ�yv$��mx�Qo�z�\k��X$��"�B\?[��Q���0ƪ��R����u��+�ݱq���Do�g9����Bӧ9�,�Kw�׾</;��xbު�y]�pK��o���o��藆ż�C����h���n���I��S�J%�;FDؒ����������b���6J,l+���O��������q�k����'@�0(J-u��_ˏ374[Ŏ⺜A�{��b����w�I1XC>��(����a,<��n�?ӝmcਨc�$��˹�B�jg2c�8�9��%3�P,N���
%`���q��\m�S���D�=�.�&&n�&2�r�S^M(���@�7i.�b�I)ޚޮ�3\C�o�E�������̇��L�d�q���=��$��y�����$�ճ���~n!�Y��_<�%G��g/����@��W����t�6V2�ˀش�؉�
HS�h��׿��vF�(�+s�=A[v4+Y������$��l�ώ z���Ø0�ӧ�>0Ԥ��+�mJ�����+�:����r��b���
w��&cU~���`+1M7��GtoΟ�D5�l�a�4�>wNk�;��䩨�(RMr�-u���k�`�q@�P^���AN`�f�5�^�Ϥ
^�fu�\q����_�W��S�h�Xn��c5�I]�iIo>hN���K��V���
���'�[�*F��U��;$��t��e���<�V�m�*Hqe�e�0�&�3"����a=�s��k��h�t\�֣��x���c�pE�:b��֊_��Zc��41��(d�z���,닲�V�|f��:�E�o�yʆV��y�Y�]̃�f�̤\�)��e�|$������^I�׭�c��:l3�3?�>�!t%Z����H�����N��I9N�� ���VL%%3�M�	���D��׶&V7$�²����
��>�)��%�|�؞ Pr�n��&�*�rwS�(��k����a'ת�aa���|�����-cJCbxt/f&#*��N&��b"C#���/��tk5�{��������7|��5��{����vDd7��.�Ӭt�h4����$��+�����.jp�Ak����%
���l��a>v���g����[vo�q�`���V|�2W��pq����8T_A��XΜh�7������lj��w�݌P����]xb�-�"R�H���_�U�{���@C>�S���P?,�+ॅ�ܘ�1���g�@�c4]�h�b?�g�,��m��WL0:Ө��2�0�54��y�?�ӷ^����v�dҽ	p��F�ԅ�A�$,�	`���y�KS�&��>���'x�/!��hW_�|���n�i��Y��~.���AZ��*#��a@B�	�A@��E�6I�Gq!(C��,Ğ&�ICx\LbI�-�){�[I�M���S�it�62��@��XӪ�� ����Àw���sQ��2�?�3,�L�!��%v�K5�g�i�����"�������D�����Pk��� US��Z��m_����ٝ�ǟBK	��v��06�=0�K!9
y�Z=�}� %�����]6���o�8Bwe���������f�"�����M9������x��E ���7�@�pM�V{�P�i��{�M�{y@�Ҽ�'ڨ��g�̶w{7e��9�ʘp���zL!"�K3�rRw'v[w{M]hT���OqH=�^�������\�2�k}ۏ�9Qs�Մ�ڒ�75��������IY�H{��E�t=ƠS�׼#X3��7�}��U�I�j�Z.�{�)Pi0�G�����c��4\Y�\�ҵ3T�۸����2:��#����\�S�.C�tv�q�ݯ�O�؜#�P-��LLs���*�<�'}D޹�f���w���z�%��_��d���W�b#�*X�h���n9��07	)Л4