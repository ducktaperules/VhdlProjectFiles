--megafunction wizard: %Altera SOPC Builder%
--GENERATION: STANDARD
--VERSION: WM1.0


--Legal Notice: (C)2011 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ad7928_spi_control_port_arbitrator is 
        port (
              -- inputs:
                 signal ad7928_spi_control_port_dataavailable : IN STD_LOGIC;
                 signal ad7928_spi_control_port_endofpacket : IN STD_LOGIC;
                 signal ad7928_spi_control_port_irq : IN STD_LOGIC;
                 signal ad7928_spi_control_port_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal ad7928_spi_control_port_readyfordata : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_2_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal gpib_edm1_clock_2_out_read : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_out_write : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal ad7928_spi_control_port_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal ad7928_spi_control_port_chipselect : OUT STD_LOGIC;
                 signal ad7928_spi_control_port_dataavailable_from_sa : OUT STD_LOGIC;
                 signal ad7928_spi_control_port_endofpacket_from_sa : OUT STD_LOGIC;
                 signal ad7928_spi_control_port_irq_from_sa : OUT STD_LOGIC;
                 signal ad7928_spi_control_port_read_n : OUT STD_LOGIC;
                 signal ad7928_spi_control_port_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal ad7928_spi_control_port_readyfordata_from_sa : OUT STD_LOGIC;
                 signal ad7928_spi_control_port_reset_n : OUT STD_LOGIC;
                 signal ad7928_spi_control_port_write_n : OUT STD_LOGIC;
                 signal ad7928_spi_control_port_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal d1_ad7928_spi_control_port_end_xfer : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_out_granted_ad7928_spi_control_port : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_out_read_data_valid_ad7928_spi_control_port : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_out_requests_ad7928_spi_control_port : OUT STD_LOGIC
              );
end entity ad7928_spi_control_port_arbitrator;


architecture europa of ad7928_spi_control_port_arbitrator is
                signal ad7928_spi_control_port_allgrants :  STD_LOGIC;
                signal ad7928_spi_control_port_allow_new_arb_cycle :  STD_LOGIC;
                signal ad7928_spi_control_port_any_bursting_master_saved_grant :  STD_LOGIC;
                signal ad7928_spi_control_port_any_continuerequest :  STD_LOGIC;
                signal ad7928_spi_control_port_arb_counter_enable :  STD_LOGIC;
                signal ad7928_spi_control_port_arb_share_counter :  STD_LOGIC;
                signal ad7928_spi_control_port_arb_share_counter_next_value :  STD_LOGIC;
                signal ad7928_spi_control_port_arb_share_set_values :  STD_LOGIC;
                signal ad7928_spi_control_port_beginbursttransfer_internal :  STD_LOGIC;
                signal ad7928_spi_control_port_begins_xfer :  STD_LOGIC;
                signal ad7928_spi_control_port_end_xfer :  STD_LOGIC;
                signal ad7928_spi_control_port_firsttransfer :  STD_LOGIC;
                signal ad7928_spi_control_port_grant_vector :  STD_LOGIC;
                signal ad7928_spi_control_port_in_a_read_cycle :  STD_LOGIC;
                signal ad7928_spi_control_port_in_a_write_cycle :  STD_LOGIC;
                signal ad7928_spi_control_port_master_qreq_vector :  STD_LOGIC;
                signal ad7928_spi_control_port_non_bursting_master_requests :  STD_LOGIC;
                signal ad7928_spi_control_port_reg_firsttransfer :  STD_LOGIC;
                signal ad7928_spi_control_port_slavearbiterlockenable :  STD_LOGIC;
                signal ad7928_spi_control_port_slavearbiterlockenable2 :  STD_LOGIC;
                signal ad7928_spi_control_port_unreg_firsttransfer :  STD_LOGIC;
                signal ad7928_spi_control_port_waits_for_read :  STD_LOGIC;
                signal ad7928_spi_control_port_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_ad7928_spi_control_port :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_arbiterlock :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_arbiterlock2 :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_continuerequest :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_saved_grant_ad7928_spi_control_port :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_gpib_edm1_clock_2_out_granted_ad7928_spi_control_port :  STD_LOGIC;
                signal internal_gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port :  STD_LOGIC;
                signal internal_gpib_edm1_clock_2_out_requests_ad7928_spi_control_port :  STD_LOGIC;
                signal wait_for_ad7928_spi_control_port_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT ad7928_spi_control_port_end_xfer;
    end if;

  end process;

  ad7928_spi_control_port_begins_xfer <= NOT d1_reasons_to_wait AND (internal_gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port);
  --assign ad7928_spi_control_port_readdata_from_sa = ad7928_spi_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  ad7928_spi_control_port_readdata_from_sa <= ad7928_spi_control_port_readdata;
  internal_gpib_edm1_clock_2_out_requests_ad7928_spi_control_port <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((gpib_edm1_clock_2_out_read OR gpib_edm1_clock_2_out_write)))))));
  --assign ad7928_spi_control_port_dataavailable_from_sa = ad7928_spi_control_port_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  ad7928_spi_control_port_dataavailable_from_sa <= ad7928_spi_control_port_dataavailable;
  --assign ad7928_spi_control_port_readyfordata_from_sa = ad7928_spi_control_port_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  ad7928_spi_control_port_readyfordata_from_sa <= ad7928_spi_control_port_readyfordata;
  --ad7928_spi_control_port_arb_share_counter set values, which is an e_mux
  ad7928_spi_control_port_arb_share_set_values <= std_logic'('1');
  --ad7928_spi_control_port_non_bursting_master_requests mux, which is an e_mux
  ad7928_spi_control_port_non_bursting_master_requests <= internal_gpib_edm1_clock_2_out_requests_ad7928_spi_control_port;
  --ad7928_spi_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  ad7928_spi_control_port_any_bursting_master_saved_grant <= std_logic'('0');
  --ad7928_spi_control_port_arb_share_counter_next_value assignment, which is an e_assign
  ad7928_spi_control_port_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(ad7928_spi_control_port_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ad7928_spi_control_port_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(ad7928_spi_control_port_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ad7928_spi_control_port_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --ad7928_spi_control_port_allgrants all slave grants, which is an e_mux
  ad7928_spi_control_port_allgrants <= ad7928_spi_control_port_grant_vector;
  --ad7928_spi_control_port_end_xfer assignment, which is an e_assign
  ad7928_spi_control_port_end_xfer <= NOT ((ad7928_spi_control_port_waits_for_read OR ad7928_spi_control_port_waits_for_write));
  --end_xfer_arb_share_counter_term_ad7928_spi_control_port arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_ad7928_spi_control_port <= ad7928_spi_control_port_end_xfer AND (((NOT ad7928_spi_control_port_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --ad7928_spi_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  ad7928_spi_control_port_arb_counter_enable <= ((end_xfer_arb_share_counter_term_ad7928_spi_control_port AND ad7928_spi_control_port_allgrants)) OR ((end_xfer_arb_share_counter_term_ad7928_spi_control_port AND NOT ad7928_spi_control_port_non_bursting_master_requests));
  --ad7928_spi_control_port_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ad7928_spi_control_port_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(ad7928_spi_control_port_arb_counter_enable) = '1' then 
        ad7928_spi_control_port_arb_share_counter <= ad7928_spi_control_port_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ad7928_spi_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ad7928_spi_control_port_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((ad7928_spi_control_port_master_qreq_vector AND end_xfer_arb_share_counter_term_ad7928_spi_control_port)) OR ((end_xfer_arb_share_counter_term_ad7928_spi_control_port AND NOT ad7928_spi_control_port_non_bursting_master_requests)))) = '1' then 
        ad7928_spi_control_port_slavearbiterlockenable <= ad7928_spi_control_port_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_2/out ad7928/spi_control_port arbiterlock, which is an e_assign
  gpib_edm1_clock_2_out_arbiterlock <= ad7928_spi_control_port_slavearbiterlockenable AND gpib_edm1_clock_2_out_continuerequest;
  --ad7928_spi_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  ad7928_spi_control_port_slavearbiterlockenable2 <= ad7928_spi_control_port_arb_share_counter_next_value;
  --gpib_edm1_clock_2/out ad7928/spi_control_port arbiterlock2, which is an e_assign
  gpib_edm1_clock_2_out_arbiterlock2 <= ad7928_spi_control_port_slavearbiterlockenable2 AND gpib_edm1_clock_2_out_continuerequest;
  --ad7928_spi_control_port_any_continuerequest at least one master continues requesting, which is an e_assign
  ad7928_spi_control_port_any_continuerequest <= std_logic'('1');
  --gpib_edm1_clock_2_out_continuerequest continued request, which is an e_assign
  gpib_edm1_clock_2_out_continuerequest <= std_logic'('1');
  internal_gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port <= internal_gpib_edm1_clock_2_out_requests_ad7928_spi_control_port;
  --ad7928_spi_control_port_writedata mux, which is an e_mux
  ad7928_spi_control_port_writedata <= gpib_edm1_clock_2_out_writedata;
  --assign ad7928_spi_control_port_endofpacket_from_sa = ad7928_spi_control_port_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  ad7928_spi_control_port_endofpacket_from_sa <= ad7928_spi_control_port_endofpacket;
  --master is always granted when requested
  internal_gpib_edm1_clock_2_out_granted_ad7928_spi_control_port <= internal_gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port;
  --gpib_edm1_clock_2/out saved-grant ad7928/spi_control_port, which is an e_assign
  gpib_edm1_clock_2_out_saved_grant_ad7928_spi_control_port <= internal_gpib_edm1_clock_2_out_requests_ad7928_spi_control_port;
  --allow new arb cycle for ad7928/spi_control_port, which is an e_assign
  ad7928_spi_control_port_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  ad7928_spi_control_port_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  ad7928_spi_control_port_master_qreq_vector <= std_logic'('1');
  --ad7928_spi_control_port_reset_n assignment, which is an e_assign
  ad7928_spi_control_port_reset_n <= reset_n;
  ad7928_spi_control_port_chipselect <= internal_gpib_edm1_clock_2_out_granted_ad7928_spi_control_port;
  --ad7928_spi_control_port_firsttransfer first transaction, which is an e_assign
  ad7928_spi_control_port_firsttransfer <= A_WE_StdLogic((std_logic'(ad7928_spi_control_port_begins_xfer) = '1'), ad7928_spi_control_port_unreg_firsttransfer, ad7928_spi_control_port_reg_firsttransfer);
  --ad7928_spi_control_port_unreg_firsttransfer first transaction, which is an e_assign
  ad7928_spi_control_port_unreg_firsttransfer <= NOT ((ad7928_spi_control_port_slavearbiterlockenable AND ad7928_spi_control_port_any_continuerequest));
  --ad7928_spi_control_port_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ad7928_spi_control_port_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(ad7928_spi_control_port_begins_xfer) = '1' then 
        ad7928_spi_control_port_reg_firsttransfer <= ad7928_spi_control_port_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --ad7928_spi_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  ad7928_spi_control_port_beginbursttransfer_internal <= ad7928_spi_control_port_begins_xfer;
  --~ad7928_spi_control_port_read_n assignment, which is an e_mux
  ad7928_spi_control_port_read_n <= NOT ((internal_gpib_edm1_clock_2_out_granted_ad7928_spi_control_port AND gpib_edm1_clock_2_out_read));
  --~ad7928_spi_control_port_write_n assignment, which is an e_mux
  ad7928_spi_control_port_write_n <= NOT ((internal_gpib_edm1_clock_2_out_granted_ad7928_spi_control_port AND gpib_edm1_clock_2_out_write));
  --ad7928_spi_control_port_address mux, which is an e_mux
  ad7928_spi_control_port_address <= gpib_edm1_clock_2_out_nativeaddress;
  --d1_ad7928_spi_control_port_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_ad7928_spi_control_port_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_ad7928_spi_control_port_end_xfer <= ad7928_spi_control_port_end_xfer;
    end if;

  end process;

  --ad7928_spi_control_port_waits_for_read in a cycle, which is an e_mux
  ad7928_spi_control_port_waits_for_read <= ad7928_spi_control_port_in_a_read_cycle AND ad7928_spi_control_port_begins_xfer;
  --ad7928_spi_control_port_in_a_read_cycle assignment, which is an e_assign
  ad7928_spi_control_port_in_a_read_cycle <= internal_gpib_edm1_clock_2_out_granted_ad7928_spi_control_port AND gpib_edm1_clock_2_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= ad7928_spi_control_port_in_a_read_cycle;
  --ad7928_spi_control_port_waits_for_write in a cycle, which is an e_mux
  ad7928_spi_control_port_waits_for_write <= ad7928_spi_control_port_in_a_write_cycle AND ad7928_spi_control_port_begins_xfer;
  --ad7928_spi_control_port_in_a_write_cycle assignment, which is an e_assign
  ad7928_spi_control_port_in_a_write_cycle <= internal_gpib_edm1_clock_2_out_granted_ad7928_spi_control_port AND gpib_edm1_clock_2_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= ad7928_spi_control_port_in_a_write_cycle;
  wait_for_ad7928_spi_control_port_counter <= std_logic'('0');
  --assign ad7928_spi_control_port_irq_from_sa = ad7928_spi_control_port_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  ad7928_spi_control_port_irq_from_sa <= ad7928_spi_control_port_irq;
  --vhdl renameroo for output signals
  gpib_edm1_clock_2_out_granted_ad7928_spi_control_port <= internal_gpib_edm1_clock_2_out_granted_ad7928_spi_control_port;
  --vhdl renameroo for output signals
  gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port <= internal_gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port;
  --vhdl renameroo for output signals
  gpib_edm1_clock_2_out_requests_ad7928_spi_control_port <= internal_gpib_edm1_clock_2_out_requests_ad7928_spi_control_port;
--synthesis translate_off
    --ad7928/spi_control_port enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_0_data_master_to_clock_crossing_0_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_0_data_master_to_clock_crossing_0_s1_module;


architecture europa of rdv_fifo_for_cpu_0_data_master_to_clock_crossing_0_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_15;
  empty <= NOT(full_0);
  full_16 <= std_logic'('0');
  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 6);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 6);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 6);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_0_instruction_master_to_clock_crossing_0_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_0_instruction_master_to_clock_crossing_0_s1_module;


architecture europa of rdv_fifo_for_cpu_0_instruction_master_to_clock_crossing_0_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_15;
  empty <= NOT(full_0);
  full_16 <= std_logic'('0');
  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 6);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 6);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 6);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity clock_crossing_0_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_s1_endofpacket : IN STD_LOGIC;
                 signal clock_crossing_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_0_s1_readdatavalid : IN STD_LOGIC;
                 signal clock_crossing_0_s1_waitrequest : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_instruction_master_read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_s1_address : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_0_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal clock_crossing_0_s1_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_s1_read : OUT STD_LOGIC;
                 signal clock_crossing_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_0_s1_reset_n : OUT STD_LOGIC;
                 signal clock_crossing_0_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal clock_crossing_0_s1_write : OUT STD_LOGIC;
                 signal clock_crossing_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_data_master_granted_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_granted_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_requests_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal d1_clock_crossing_0_s1_end_xfer : OUT STD_LOGIC
              );
end entity clock_crossing_0_s1_arbitrator;


architecture europa of clock_crossing_0_s1_arbitrator is
component rdv_fifo_for_cpu_0_data_master_to_clock_crossing_0_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_0_data_master_to_clock_crossing_0_s1_module;

component rdv_fifo_for_cpu_0_instruction_master_to_clock_crossing_0_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_0_instruction_master_to_clock_crossing_0_s1_module;

                signal clock_crossing_0_s1_allgrants :  STD_LOGIC;
                signal clock_crossing_0_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal clock_crossing_0_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal clock_crossing_0_s1_any_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal clock_crossing_0_s1_arb_counter_enable :  STD_LOGIC;
                signal clock_crossing_0_s1_arb_share_counter :  STD_LOGIC;
                signal clock_crossing_0_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal clock_crossing_0_s1_arb_share_set_values :  STD_LOGIC;
                signal clock_crossing_0_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal clock_crossing_0_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal clock_crossing_0_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal clock_crossing_0_s1_begins_xfer :  STD_LOGIC;
                signal clock_crossing_0_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clock_crossing_0_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal clock_crossing_0_s1_end_xfer :  STD_LOGIC;
                signal clock_crossing_0_s1_firsttransfer :  STD_LOGIC;
                signal clock_crossing_0_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal clock_crossing_0_s1_in_a_read_cycle :  STD_LOGIC;
                signal clock_crossing_0_s1_in_a_write_cycle :  STD_LOGIC;
                signal clock_crossing_0_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal clock_crossing_0_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal clock_crossing_0_s1_non_bursting_master_requests :  STD_LOGIC;
                signal clock_crossing_0_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal clock_crossing_0_s1_reg_firsttransfer :  STD_LOGIC;
                signal clock_crossing_0_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal clock_crossing_0_s1_slavearbiterlockenable :  STD_LOGIC;
                signal clock_crossing_0_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal clock_crossing_0_s1_unreg_firsttransfer :  STD_LOGIC;
                signal clock_crossing_0_s1_waits_for_read :  STD_LOGIC;
                signal clock_crossing_0_s1_waits_for_write :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_rdv_fifo_empty_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_data_master_rdv_fifo_output_from_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_0_instruction_master_rdv_fifo_empty_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_rdv_fifo_output_from_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_saved_grant_clock_crossing_0_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_clock_crossing_0_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_s1_waitrequest_from_sa :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_clock_crossing_0_s1 :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_clock_crossing_0_s1 :  STD_LOGIC;
                signal internal_cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_clock_crossing_0_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_granted_clock_crossing_0_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_requests_clock_crossing_0_s1 :  STD_LOGIC;
                signal last_cycle_cpu_0_data_master_granted_slave_clock_crossing_0_s1 :  STD_LOGIC;
                signal last_cycle_cpu_0_instruction_master_granted_slave_clock_crossing_0_s1 :  STD_LOGIC;
                signal module_input :  STD_LOGIC;
                signal module_input1 :  STD_LOGIC;
                signal module_input2 :  STD_LOGIC;
                signal module_input3 :  STD_LOGIC;
                signal module_input4 :  STD_LOGIC;
                signal module_input5 :  STD_LOGIC;
                signal shifted_address_to_clock_crossing_0_s1_from_cpu_0_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal shifted_address_to_clock_crossing_0_s1_from_cpu_0_instruction_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_clock_crossing_0_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT clock_crossing_0_s1_end_xfer;
    end if;

  end process;

  clock_crossing_0_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpu_0_data_master_qualified_request_clock_crossing_0_s1 OR internal_cpu_0_instruction_master_qualified_request_clock_crossing_0_s1));
  --assign clock_crossing_0_s1_readdata_from_sa = clock_crossing_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  clock_crossing_0_s1_readdata_from_sa <= clock_crossing_0_s1_readdata;
  internal_cpu_0_data_master_requests_clock_crossing_0_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(27 DOWNTO 8) & std_logic_vector'("00000000")) = std_logic_vector'("1001000000000000000000000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign clock_crossing_0_s1_waitrequest_from_sa = clock_crossing_0_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_clock_crossing_0_s1_waitrequest_from_sa <= clock_crossing_0_s1_waitrequest;
  --assign clock_crossing_0_s1_readdatavalid_from_sa = clock_crossing_0_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  clock_crossing_0_s1_readdatavalid_from_sa <= clock_crossing_0_s1_readdatavalid;
  --clock_crossing_0_s1_arb_share_counter set values, which is an e_mux
  clock_crossing_0_s1_arb_share_set_values <= std_logic'('1');
  --clock_crossing_0_s1_non_bursting_master_requests mux, which is an e_mux
  clock_crossing_0_s1_non_bursting_master_requests <= ((internal_cpu_0_data_master_requests_clock_crossing_0_s1 OR internal_cpu_0_instruction_master_requests_clock_crossing_0_s1) OR internal_cpu_0_data_master_requests_clock_crossing_0_s1) OR internal_cpu_0_instruction_master_requests_clock_crossing_0_s1;
  --clock_crossing_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  clock_crossing_0_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --clock_crossing_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  clock_crossing_0_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(clock_crossing_0_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(clock_crossing_0_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --clock_crossing_0_s1_allgrants all slave grants, which is an e_mux
  clock_crossing_0_s1_allgrants <= (((or_reduce(clock_crossing_0_s1_grant_vector)) OR (or_reduce(clock_crossing_0_s1_grant_vector))) OR (or_reduce(clock_crossing_0_s1_grant_vector))) OR (or_reduce(clock_crossing_0_s1_grant_vector));
  --clock_crossing_0_s1_end_xfer assignment, which is an e_assign
  clock_crossing_0_s1_end_xfer <= NOT ((clock_crossing_0_s1_waits_for_read OR clock_crossing_0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_clock_crossing_0_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_clock_crossing_0_s1 <= clock_crossing_0_s1_end_xfer AND (((NOT clock_crossing_0_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --clock_crossing_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  clock_crossing_0_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_clock_crossing_0_s1 AND clock_crossing_0_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_clock_crossing_0_s1 AND NOT clock_crossing_0_s1_non_bursting_master_requests));
  --clock_crossing_0_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_0_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(clock_crossing_0_s1_arb_counter_enable) = '1' then 
        clock_crossing_0_s1_arb_share_counter <= clock_crossing_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_0_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(clock_crossing_0_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_clock_crossing_0_s1)) OR ((end_xfer_arb_share_counter_term_clock_crossing_0_s1 AND NOT clock_crossing_0_s1_non_bursting_master_requests)))) = '1' then 
        clock_crossing_0_s1_slavearbiterlockenable <= clock_crossing_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_0/data_master clock_crossing_0/s1 arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= clock_crossing_0_s1_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --clock_crossing_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  clock_crossing_0_s1_slavearbiterlockenable2 <= clock_crossing_0_s1_arb_share_counter_next_value;
  --cpu_0/data_master clock_crossing_0/s1 arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= clock_crossing_0_s1_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --cpu_0/instruction_master clock_crossing_0/s1 arbiterlock, which is an e_assign
  cpu_0_instruction_master_arbiterlock <= clock_crossing_0_s1_slavearbiterlockenable AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master clock_crossing_0/s1 arbiterlock2, which is an e_assign
  cpu_0_instruction_master_arbiterlock2 <= clock_crossing_0_s1_slavearbiterlockenable2 AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master granted clock_crossing_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_instruction_master_granted_slave_clock_crossing_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_instruction_master_granted_slave_clock_crossing_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_instruction_master_saved_grant_clock_crossing_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((clock_crossing_0_s1_arbitration_holdoff_internal OR NOT internal_cpu_0_instruction_master_requests_clock_crossing_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_instruction_master_granted_slave_clock_crossing_0_s1))))));
    end if;

  end process;

  --cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  cpu_0_instruction_master_continuerequest <= last_cycle_cpu_0_instruction_master_granted_slave_clock_crossing_0_s1 AND internal_cpu_0_instruction_master_requests_clock_crossing_0_s1;
  --clock_crossing_0_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  clock_crossing_0_s1_any_continuerequest <= cpu_0_instruction_master_continuerequest OR cpu_0_data_master_continuerequest;
  internal_cpu_0_data_master_qualified_request_clock_crossing_0_s1 <= internal_cpu_0_data_master_requests_clock_crossing_0_s1 AND NOT (((((cpu_0_data_master_read AND ((NOT cpu_0_data_master_waitrequest OR (internal_cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register))))) OR (((NOT cpu_0_data_master_waitrequest) AND cpu_0_data_master_write))) OR cpu_0_instruction_master_arbiterlock));
  --unique name for clock_crossing_0_s1_move_on_to_next_transaction, which is an e_assign
  clock_crossing_0_s1_move_on_to_next_transaction <= clock_crossing_0_s1_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_0_data_master_to_clock_crossing_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_0_data_master_to_clock_crossing_0_s1 : rdv_fifo_for_cpu_0_data_master_to_clock_crossing_0_s1_module
    port map(
      data_out => cpu_0_data_master_rdv_fifo_output_from_clock_crossing_0_s1,
      empty => open,
      fifo_contains_ones_n => cpu_0_data_master_rdv_fifo_empty_clock_crossing_0_s1,
      full => open,
      clear_fifo => module_input,
      clk => clk,
      data_in => internal_cpu_0_data_master_granted_clock_crossing_0_s1,
      read => clock_crossing_0_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input1,
      write => module_input2
    );

  module_input <= std_logic'('0');
  module_input1 <= std_logic'('0');
  module_input2 <= in_a_read_cycle AND NOT clock_crossing_0_s1_waits_for_read;

  internal_cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register <= NOT cpu_0_data_master_rdv_fifo_empty_clock_crossing_0_s1;
  --local readdatavalid cpu_0_data_master_read_data_valid_clock_crossing_0_s1, which is an e_mux
  cpu_0_data_master_read_data_valid_clock_crossing_0_s1 <= ((clock_crossing_0_s1_readdatavalid_from_sa AND cpu_0_data_master_rdv_fifo_output_from_clock_crossing_0_s1)) AND NOT cpu_0_data_master_rdv_fifo_empty_clock_crossing_0_s1;
  --clock_crossing_0_s1_writedata mux, which is an e_mux
  clock_crossing_0_s1_writedata <= cpu_0_data_master_writedata;
  --assign clock_crossing_0_s1_endofpacket_from_sa = clock_crossing_0_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  clock_crossing_0_s1_endofpacket_from_sa <= clock_crossing_0_s1_endofpacket;
  internal_cpu_0_instruction_master_requests_clock_crossing_0_s1 <= ((to_std_logic(((Std_Logic_Vector'(cpu_0_instruction_master_address_to_slave(27 DOWNTO 8) & std_logic_vector'("00000000")) = std_logic_vector'("1001000000000000000000000000")))) AND (cpu_0_instruction_master_read))) AND cpu_0_instruction_master_read;
  --cpu_0/data_master granted clock_crossing_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_data_master_granted_slave_clock_crossing_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_data_master_granted_slave_clock_crossing_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_data_master_saved_grant_clock_crossing_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((clock_crossing_0_s1_arbitration_holdoff_internal OR NOT internal_cpu_0_data_master_requests_clock_crossing_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_data_master_granted_slave_clock_crossing_0_s1))))));
    end if;

  end process;

  --cpu_0_data_master_continuerequest continued request, which is an e_mux
  cpu_0_data_master_continuerequest <= last_cycle_cpu_0_data_master_granted_slave_clock_crossing_0_s1 AND internal_cpu_0_data_master_requests_clock_crossing_0_s1;
  internal_cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 <= internal_cpu_0_instruction_master_requests_clock_crossing_0_s1 AND NOT ((((cpu_0_instruction_master_read AND (internal_cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register))) OR cpu_0_data_master_arbiterlock));
  --rdv_fifo_for_cpu_0_instruction_master_to_clock_crossing_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_0_instruction_master_to_clock_crossing_0_s1 : rdv_fifo_for_cpu_0_instruction_master_to_clock_crossing_0_s1_module
    port map(
      data_out => cpu_0_instruction_master_rdv_fifo_output_from_clock_crossing_0_s1,
      empty => open,
      fifo_contains_ones_n => cpu_0_instruction_master_rdv_fifo_empty_clock_crossing_0_s1,
      full => open,
      clear_fifo => module_input3,
      clk => clk,
      data_in => internal_cpu_0_instruction_master_granted_clock_crossing_0_s1,
      read => clock_crossing_0_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input4,
      write => module_input5
    );

  module_input3 <= std_logic'('0');
  module_input4 <= std_logic'('0');
  module_input5 <= in_a_read_cycle AND NOT clock_crossing_0_s1_waits_for_read;

  internal_cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register <= NOT cpu_0_instruction_master_rdv_fifo_empty_clock_crossing_0_s1;
  --local readdatavalid cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1, which is an e_mux
  cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1 <= ((clock_crossing_0_s1_readdatavalid_from_sa AND cpu_0_instruction_master_rdv_fifo_output_from_clock_crossing_0_s1)) AND NOT cpu_0_instruction_master_rdv_fifo_empty_clock_crossing_0_s1;
  --allow new arb cycle for clock_crossing_0/s1, which is an e_assign
  clock_crossing_0_s1_allow_new_arb_cycle <= NOT cpu_0_data_master_arbiterlock AND NOT cpu_0_instruction_master_arbiterlock;
  --cpu_0/instruction_master assignment into master qualified-requests vector for clock_crossing_0/s1, which is an e_assign
  clock_crossing_0_s1_master_qreq_vector(0) <= internal_cpu_0_instruction_master_qualified_request_clock_crossing_0_s1;
  --cpu_0/instruction_master grant clock_crossing_0/s1, which is an e_assign
  internal_cpu_0_instruction_master_granted_clock_crossing_0_s1 <= clock_crossing_0_s1_grant_vector(0);
  --cpu_0/instruction_master saved-grant clock_crossing_0/s1, which is an e_assign
  cpu_0_instruction_master_saved_grant_clock_crossing_0_s1 <= clock_crossing_0_s1_arb_winner(0) AND internal_cpu_0_instruction_master_requests_clock_crossing_0_s1;
  --cpu_0/data_master assignment into master qualified-requests vector for clock_crossing_0/s1, which is an e_assign
  clock_crossing_0_s1_master_qreq_vector(1) <= internal_cpu_0_data_master_qualified_request_clock_crossing_0_s1;
  --cpu_0/data_master grant clock_crossing_0/s1, which is an e_assign
  internal_cpu_0_data_master_granted_clock_crossing_0_s1 <= clock_crossing_0_s1_grant_vector(1);
  --cpu_0/data_master saved-grant clock_crossing_0/s1, which is an e_assign
  cpu_0_data_master_saved_grant_clock_crossing_0_s1 <= clock_crossing_0_s1_arb_winner(1) AND internal_cpu_0_data_master_requests_clock_crossing_0_s1;
  --clock_crossing_0/s1 chosen-master double-vector, which is an e_assign
  clock_crossing_0_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((clock_crossing_0_s1_master_qreq_vector & clock_crossing_0_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT clock_crossing_0_s1_master_qreq_vector & NOT clock_crossing_0_s1_master_qreq_vector))) + (std_logic_vector'("000") & (clock_crossing_0_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  clock_crossing_0_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((clock_crossing_0_s1_allow_new_arb_cycle AND or_reduce(clock_crossing_0_s1_grant_vector)))) = '1'), clock_crossing_0_s1_grant_vector, clock_crossing_0_s1_saved_chosen_master_vector);
  --saved clock_crossing_0_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_0_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(clock_crossing_0_s1_allow_new_arb_cycle) = '1' then 
        clock_crossing_0_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(clock_crossing_0_s1_grant_vector)) = '1'), clock_crossing_0_s1_grant_vector, clock_crossing_0_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  clock_crossing_0_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((clock_crossing_0_s1_chosen_master_double_vector(1) OR clock_crossing_0_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((clock_crossing_0_s1_chosen_master_double_vector(0) OR clock_crossing_0_s1_chosen_master_double_vector(2)))));
  --clock_crossing_0/s1 chosen master rotated left, which is an e_assign
  clock_crossing_0_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(clock_crossing_0_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(clock_crossing_0_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --clock_crossing_0/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_0_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(clock_crossing_0_s1_grant_vector)) = '1' then 
        clock_crossing_0_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(clock_crossing_0_s1_end_xfer) = '1'), clock_crossing_0_s1_chosen_master_rot_left, clock_crossing_0_s1_grant_vector);
      end if;
    end if;

  end process;

  --clock_crossing_0_s1_reset_n assignment, which is an e_assign
  clock_crossing_0_s1_reset_n <= reset_n;
  --clock_crossing_0_s1_firsttransfer first transaction, which is an e_assign
  clock_crossing_0_s1_firsttransfer <= A_WE_StdLogic((std_logic'(clock_crossing_0_s1_begins_xfer) = '1'), clock_crossing_0_s1_unreg_firsttransfer, clock_crossing_0_s1_reg_firsttransfer);
  --clock_crossing_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  clock_crossing_0_s1_unreg_firsttransfer <= NOT ((clock_crossing_0_s1_slavearbiterlockenable AND clock_crossing_0_s1_any_continuerequest));
  --clock_crossing_0_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_0_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(clock_crossing_0_s1_begins_xfer) = '1' then 
        clock_crossing_0_s1_reg_firsttransfer <= clock_crossing_0_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --clock_crossing_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  clock_crossing_0_s1_beginbursttransfer_internal <= clock_crossing_0_s1_begins_xfer;
  --clock_crossing_0_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  clock_crossing_0_s1_arbitration_holdoff_internal <= clock_crossing_0_s1_begins_xfer AND clock_crossing_0_s1_firsttransfer;
  --clock_crossing_0_s1_read assignment, which is an e_mux
  clock_crossing_0_s1_read <= ((internal_cpu_0_data_master_granted_clock_crossing_0_s1 AND cpu_0_data_master_read)) OR ((internal_cpu_0_instruction_master_granted_clock_crossing_0_s1 AND cpu_0_instruction_master_read));
  --clock_crossing_0_s1_write assignment, which is an e_mux
  clock_crossing_0_s1_write <= internal_cpu_0_data_master_granted_clock_crossing_0_s1 AND cpu_0_data_master_write;
  shifted_address_to_clock_crossing_0_s1_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --clock_crossing_0_s1_address mux, which is an e_mux
  clock_crossing_0_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_clock_crossing_0_s1)) = '1'), (A_SRL(shifted_address_to_clock_crossing_0_s1_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_clock_crossing_0_s1_from_cpu_0_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 6);
  shifted_address_to_clock_crossing_0_s1_from_cpu_0_instruction_master <= cpu_0_instruction_master_address_to_slave;
  --slaveid clock_crossing_0_s1_nativeaddress nativeaddress mux, which is an e_mux
  clock_crossing_0_s1_nativeaddress <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_clock_crossing_0_s1)) = '1'), (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(cpu_0_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")))), 6);
  --d1_clock_crossing_0_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_clock_crossing_0_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_clock_crossing_0_s1_end_xfer <= clock_crossing_0_s1_end_xfer;
    end if;

  end process;

  --clock_crossing_0_s1_waits_for_read in a cycle, which is an e_mux
  clock_crossing_0_s1_waits_for_read <= clock_crossing_0_s1_in_a_read_cycle AND internal_clock_crossing_0_s1_waitrequest_from_sa;
  --clock_crossing_0_s1_in_a_read_cycle assignment, which is an e_assign
  clock_crossing_0_s1_in_a_read_cycle <= ((internal_cpu_0_data_master_granted_clock_crossing_0_s1 AND cpu_0_data_master_read)) OR ((internal_cpu_0_instruction_master_granted_clock_crossing_0_s1 AND cpu_0_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= clock_crossing_0_s1_in_a_read_cycle;
  --clock_crossing_0_s1_waits_for_write in a cycle, which is an e_mux
  clock_crossing_0_s1_waits_for_write <= clock_crossing_0_s1_in_a_write_cycle AND internal_clock_crossing_0_s1_waitrequest_from_sa;
  --clock_crossing_0_s1_in_a_write_cycle assignment, which is an e_assign
  clock_crossing_0_s1_in_a_write_cycle <= internal_cpu_0_data_master_granted_clock_crossing_0_s1 AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= clock_crossing_0_s1_in_a_write_cycle;
  wait_for_clock_crossing_0_s1_counter <= std_logic'('0');
  --clock_crossing_0_s1_byteenable byte enable port mux, which is an e_mux
  clock_crossing_0_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_clock_crossing_0_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  clock_crossing_0_s1_waitrequest_from_sa <= internal_clock_crossing_0_s1_waitrequest_from_sa;
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_clock_crossing_0_s1 <= internal_cpu_0_data_master_granted_clock_crossing_0_s1;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_clock_crossing_0_s1 <= internal_cpu_0_data_master_qualified_request_clock_crossing_0_s1;
  --vhdl renameroo for output signals
  cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register <= internal_cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_clock_crossing_0_s1 <= internal_cpu_0_data_master_requests_clock_crossing_0_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_granted_clock_crossing_0_s1 <= internal_cpu_0_instruction_master_granted_clock_crossing_0_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 <= internal_cpu_0_instruction_master_qualified_request_clock_crossing_0_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register <= internal_cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_requests_clock_crossing_0_s1 <= internal_cpu_0_instruction_master_requests_clock_crossing_0_s1;
--synthesis translate_off
    --clock_crossing_0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_data_master_granted_clock_crossing_0_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_instruction_master_granted_clock_crossing_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line, now);
          write(write_line, string'(": "));
          write(write_line, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line.all);
          deallocate (write_line);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line1 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_saved_grant_clock_crossing_0_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_saved_grant_clock_crossing_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line1, now);
          write(write_line1, string'(": "));
          write(write_line1, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line1.all);
          deallocate (write_line1);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity clock_crossing_0_m1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_0_m1_granted_gpib_edm1_clock_2_in : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_gpib_edm1_clock_3_in : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_gpib_leds_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_gpio1_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_gpio2_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_high_res_timer_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_led_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_sys_clk_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_gpib_leds_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_gpio1_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_gpio2_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_high_res_timer_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_led_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_sys_clk_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_gpib_leds_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_gpio1_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_gpio2_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_high_res_timer_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_led_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_sys_clk_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_gpib_edm1_clock_2_in : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_gpib_edm1_clock_3_in : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_gpib_leds_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_gpio1_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_gpio2_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_high_res_timer_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_led_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_sys_clk_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_gpib_edm1_clock_2_in_end_xfer : IN STD_LOGIC;
                 signal d1_gpib_edm1_clock_3_in_end_xfer : IN STD_LOGIC;
                 signal d1_gpib_leds_s1_end_xfer : IN STD_LOGIC;
                 signal d1_gpio1_s1_end_xfer : IN STD_LOGIC;
                 signal d1_gpio2_s1_end_xfer : IN STD_LOGIC;
                 signal d1_high_res_timer_s1_end_xfer : IN STD_LOGIC;
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                 signal d1_led_pio_s1_end_xfer : IN STD_LOGIC;
                 signal d1_sys_clk_s1_end_xfer : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_in_endofpacket_from_sa : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_2_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_in_endofpacket_from_sa : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_3_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal gpib_leds_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gpio1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gpio2_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal high_res_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal led_pio_s1_readdata_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal clock_crossing_0_m1_address_to_slave : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_endofpacket : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_latency_counter : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_0_m1_readdatavalid : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_reset_n : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_waitrequest : OUT STD_LOGIC
              );
end entity clock_crossing_0_m1_arbitrator;


architecture europa of clock_crossing_0_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal clock_crossing_0_m1_address_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal clock_crossing_0_m1_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clock_crossing_0_m1_is_granted_some_slave :  STD_LOGIC;
                signal clock_crossing_0_m1_read_but_no_slave_selected :  STD_LOGIC;
                signal clock_crossing_0_m1_read_last_time :  STD_LOGIC;
                signal clock_crossing_0_m1_run :  STD_LOGIC;
                signal clock_crossing_0_m1_write_last_time :  STD_LOGIC;
                signal clock_crossing_0_m1_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_clock_crossing_0_m1_address_to_slave :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_clock_crossing_0_m1_latency_counter :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_clock_crossing_0_m1_latency_counter :  STD_LOGIC;
                signal pre_flush_clock_crossing_0_m1_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in OR NOT clock_crossing_0_m1_requests_gpib_edm1_clock_2_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in OR NOT ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT gpib_edm1_clock_2_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in OR NOT ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT gpib_edm1_clock_2_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in OR NOT clock_crossing_0_m1_requests_gpib_edm1_clock_3_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in OR NOT ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT gpib_edm1_clock_3_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in OR NOT ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT gpib_edm1_clock_3_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_gpib_leds_s1 OR NOT clock_crossing_0_m1_requests_gpib_leds_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_gpib_leds_s1 OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_gpib_leds_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_gpib_leds_s1 OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_gpio1_s1 OR NOT clock_crossing_0_m1_requests_gpio1_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_gpio1_s1 OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_gpio1_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_gpio1_s1 OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_gpio2_s1 OR NOT clock_crossing_0_m1_requests_gpio2_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_gpio2_s1 OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_gpio2_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_gpio2_s1 OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))));
  --cascaded wait assignment, which is an e_assign
  clock_crossing_0_m1_run <= r_1 AND r_2;
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_high_res_timer_s1 OR NOT clock_crossing_0_m1_requests_high_res_timer_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_high_res_timer_s1 OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_high_res_timer_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_high_res_timer_s1 OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave OR NOT clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave OR NOT ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave OR NOT ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_led_pio_s1 OR NOT clock_crossing_0_m1_requests_led_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_led_pio_s1 OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_led_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_led_pio_s1 OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_sys_clk_s1 OR NOT clock_crossing_0_m1_requests_sys_clk_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_sys_clk_s1 OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sys_clk_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_sys_clk_s1 OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_clock_crossing_0_m1_address_to_slave <= clock_crossing_0_m1_address(7 DOWNTO 0);
  --clock_crossing_0_m1_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_0_m1_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      clock_crossing_0_m1_read_but_no_slave_selected <= (clock_crossing_0_m1_read AND clock_crossing_0_m1_run) AND NOT clock_crossing_0_m1_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  clock_crossing_0_m1_is_granted_some_slave <= (((((((clock_crossing_0_m1_granted_gpib_edm1_clock_2_in OR clock_crossing_0_m1_granted_gpib_edm1_clock_3_in) OR clock_crossing_0_m1_granted_gpib_leds_s1) OR clock_crossing_0_m1_granted_gpio1_s1) OR clock_crossing_0_m1_granted_gpio2_s1) OR clock_crossing_0_m1_granted_high_res_timer_s1) OR clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave) OR clock_crossing_0_m1_granted_led_pio_s1) OR clock_crossing_0_m1_granted_sys_clk_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_clock_crossing_0_m1_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  clock_crossing_0_m1_readdatavalid <= (((((((((((((((((((((((((clock_crossing_0_m1_read_but_no_slave_selected OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_gpib_leds_s1) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_gpio1_s1) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_gpio2_s1) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_high_res_timer_s1) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_led_pio_s1) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_sys_clk_s1;
  --clock_crossing_0/m1 readdata mux, which is an e_mux
  clock_crossing_0_m1_readdata <= (((((((((A_REP(NOT ((clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("0000000000000000") & (gpib_edm1_clock_2_in_readdata_from_sa)))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("0000000000000000") & (gpib_edm1_clock_3_in_readdata_from_sa))))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_gpib_leds_s1 AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (gpib_leds_s1_readdata_from_sa))))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_gpio1_s1 AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (gpio1_s1_readdata_from_sa))))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_gpio2_s1 AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (gpio2_s1_readdata_from_sa))))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_high_res_timer_s1 AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("0000000000000000") & (high_res_timer_s1_readdata_from_sa))))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave AND clock_crossing_0_m1_read)) , 32) OR jtag_uart_avalon_jtag_slave_readdata_from_sa))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_led_pio_s1 AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_pio_s1_readdata_from_sa)))))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_sys_clk_s1 AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("0000000000000000") & (sys_clk_s1_readdata_from_sa))));
  --actual waitrequest port, which is an e_assign
  internal_clock_crossing_0_m1_waitrequest <= NOT clock_crossing_0_m1_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_clock_crossing_0_m1_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_clock_crossing_0_m1_latency_counter <= p1_clock_crossing_0_m1_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_clock_crossing_0_m1_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((clock_crossing_0_m1_run AND clock_crossing_0_m1_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_clock_crossing_0_m1_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_clock_crossing_0_m1_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --clock_crossing_0_m1_reset_n assignment, which is an e_assign
  clock_crossing_0_m1_reset_n <= reset_n;
  --mux clock_crossing_0_m1_endofpacket, which is an e_mux
  clock_crossing_0_m1_endofpacket <= A_WE_StdLogic((std_logic'((clock_crossing_0_m1_requests_gpib_edm1_clock_2_in)) = '1'), gpib_edm1_clock_2_in_endofpacket_from_sa, gpib_edm1_clock_3_in_endofpacket_from_sa);
  --vhdl renameroo for output signals
  clock_crossing_0_m1_address_to_slave <= internal_clock_crossing_0_m1_address_to_slave;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_latency_counter <= internal_clock_crossing_0_m1_latency_counter;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_waitrequest <= internal_clock_crossing_0_m1_waitrequest;
--synthesis translate_off
    --clock_crossing_0_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_0_m1_address_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        clock_crossing_0_m1_address_last_time <= clock_crossing_0_m1_address;
      end if;

    end process;

    --clock_crossing_0/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_clock_crossing_0_m1_waitrequest AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
      end if;

    end process;

    --clock_crossing_0_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line2 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((clock_crossing_0_m1_address /= clock_crossing_0_m1_address_last_time))))) = '1' then 
          write(write_line2, now);
          write(write_line2, string'(": "));
          write(write_line2, string'("clock_crossing_0_m1_address did not heed wait!!!"));
          write(output, write_line2.all);
          deallocate (write_line2);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_0_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_0_m1_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        clock_crossing_0_m1_byteenable_last_time <= clock_crossing_0_m1_byteenable;
      end if;

    end process;

    --clock_crossing_0_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line3 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((clock_crossing_0_m1_byteenable /= clock_crossing_0_m1_byteenable_last_time))))) = '1' then 
          write(write_line3, now);
          write(write_line3, string'(": "));
          write(write_line3, string'("clock_crossing_0_m1_byteenable did not heed wait!!!"));
          write(output, write_line3.all);
          deallocate (write_line3);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_0_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_0_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        clock_crossing_0_m1_read_last_time <= clock_crossing_0_m1_read;
      end if;

    end process;

    --clock_crossing_0_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line4 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(clock_crossing_0_m1_read) /= std_logic'(clock_crossing_0_m1_read_last_time)))))) = '1' then 
          write(write_line4, now);
          write(write_line4, string'(": "));
          write(write_line4, string'("clock_crossing_0_m1_read did not heed wait!!!"));
          write(output, write_line4.all);
          deallocate (write_line4);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_0_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_0_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        clock_crossing_0_m1_write_last_time <= clock_crossing_0_m1_write;
      end if;

    end process;

    --clock_crossing_0_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line5 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(clock_crossing_0_m1_write) /= std_logic'(clock_crossing_0_m1_write_last_time)))))) = '1' then 
          write(write_line5, now);
          write(write_line5, string'(": "));
          write(write_line5, string'("clock_crossing_0_m1_write did not heed wait!!!"));
          write(output, write_line5.all);
          deallocate (write_line5);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_0_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_0_m1_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        clock_crossing_0_m1_writedata_last_time <= clock_crossing_0_m1_writedata;
      end if;

    end process;

    --clock_crossing_0_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line6 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((clock_crossing_0_m1_writedata /= clock_crossing_0_m1_writedata_last_time)))) AND clock_crossing_0_m1_write)) = '1' then 
          write(write_line6, now);
          write(write_line6, string'(": "));
          write(write_line6, string'("clock_crossing_0_m1_writedata did not heed wait!!!"));
          write(output, write_line6.all);
          deallocate (write_line6);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity clock_crossing_0_bridge_arbitrator is 
end entity clock_crossing_0_bridge_arbitrator;


architecture europa of clock_crossing_0_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_0_jtag_debug_module_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_instruction_master_read : IN STD_LOGIC;
                 signal cpu_0_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_jtag_debug_module_resetrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_granted_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_requests_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal cpu_0_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_jtag_debug_module_chipselect : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_jtag_debug_module_reset_n : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_write : OUT STD_LOGIC;
                 signal cpu_0_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_0_jtag_debug_module_end_xfer : OUT STD_LOGIC
              );
end entity cpu_0_jtag_debug_module_arbitrator;


architecture europa of cpu_0_jtag_debug_module_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_allgrants :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_allow_new_arb_cycle :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_any_continuerequest :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_arb_counter_enable :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_arb_share_counter :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_arb_share_counter_next_value :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_arb_share_set_values :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_arbitration_holdoff_internal :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_beginbursttransfer_internal :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_begins_xfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_0_jtag_debug_module_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_firsttransfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_in_a_read_cycle :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_in_a_write_cycle :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_non_bursting_master_requests :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_reg_firsttransfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_0_jtag_debug_module_slavearbiterlockenable :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_slavearbiterlockenable2 :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_unreg_firsttransfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_waits_for_read :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_cpu_0_jtag_debug_module_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cpu_0_jtag_debug_module_end_xfer;
    end if;

  end process;

  cpu_0_jtag_debug_module_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module OR internal_cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module));
  --assign cpu_0_jtag_debug_module_readdata_from_sa = cpu_0_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_0_jtag_debug_module_readdata_from_sa <= cpu_0_jtag_debug_module_readdata;
  internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(27 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("1010000000001000100000000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --cpu_0_jtag_debug_module_arb_share_counter set values, which is an e_mux
  cpu_0_jtag_debug_module_arb_share_set_values <= std_logic'('1');
  --cpu_0_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  cpu_0_jtag_debug_module_non_bursting_master_requests <= ((internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module OR internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module) OR internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module) OR internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  --cpu_0_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  cpu_0_jtag_debug_module_any_bursting_master_saved_grant <= std_logic'('0');
  --cpu_0_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  cpu_0_jtag_debug_module_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_jtag_debug_module_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_jtag_debug_module_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(cpu_0_jtag_debug_module_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_jtag_debug_module_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --cpu_0_jtag_debug_module_allgrants all slave grants, which is an e_mux
  cpu_0_jtag_debug_module_allgrants <= (((or_reduce(cpu_0_jtag_debug_module_grant_vector)) OR (or_reduce(cpu_0_jtag_debug_module_grant_vector))) OR (or_reduce(cpu_0_jtag_debug_module_grant_vector))) OR (or_reduce(cpu_0_jtag_debug_module_grant_vector));
  --cpu_0_jtag_debug_module_end_xfer assignment, which is an e_assign
  cpu_0_jtag_debug_module_end_xfer <= NOT ((cpu_0_jtag_debug_module_waits_for_read OR cpu_0_jtag_debug_module_waits_for_write));
  --end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module <= cpu_0_jtag_debug_module_end_xfer AND (((NOT cpu_0_jtag_debug_module_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cpu_0_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  cpu_0_jtag_debug_module_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module AND cpu_0_jtag_debug_module_allgrants)) OR ((end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module AND NOT cpu_0_jtag_debug_module_non_bursting_master_requests));
  --cpu_0_jtag_debug_module_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_jtag_debug_module_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_0_jtag_debug_module_arb_counter_enable) = '1' then 
        cpu_0_jtag_debug_module_arb_share_counter <= cpu_0_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_0_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_jtag_debug_module_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(cpu_0_jtag_debug_module_master_qreq_vector) AND end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module)) OR ((end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module AND NOT cpu_0_jtag_debug_module_non_bursting_master_requests)))) = '1' then 
        cpu_0_jtag_debug_module_slavearbiterlockenable <= cpu_0_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_0/data_master cpu_0/jtag_debug_module arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= cpu_0_jtag_debug_module_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --cpu_0_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cpu_0_jtag_debug_module_slavearbiterlockenable2 <= cpu_0_jtag_debug_module_arb_share_counter_next_value;
  --cpu_0/data_master cpu_0/jtag_debug_module arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= cpu_0_jtag_debug_module_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --cpu_0/instruction_master cpu_0/jtag_debug_module arbiterlock, which is an e_assign
  cpu_0_instruction_master_arbiterlock <= cpu_0_jtag_debug_module_slavearbiterlockenable AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master cpu_0/jtag_debug_module arbiterlock2, which is an e_assign
  cpu_0_instruction_master_arbiterlock2 <= cpu_0_jtag_debug_module_slavearbiterlockenable2 AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master granted cpu_0/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpu_0_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module))))));
    end if;

  end process;

  --cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  cpu_0_instruction_master_continuerequest <= last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module AND internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  --cpu_0_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  cpu_0_jtag_debug_module_any_continuerequest <= cpu_0_instruction_master_continuerequest OR cpu_0_data_master_continuerequest;
  internal_cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module <= internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module AND NOT (((((NOT cpu_0_data_master_waitrequest) AND cpu_0_data_master_write)) OR cpu_0_instruction_master_arbiterlock));
  --cpu_0_jtag_debug_module_writedata mux, which is an e_mux
  cpu_0_jtag_debug_module_writedata <= cpu_0_data_master_writedata;
  internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module <= ((to_std_logic(((Std_Logic_Vector'(cpu_0_instruction_master_address_to_slave(27 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("1010000000001000100000000000")))) AND (cpu_0_instruction_master_read))) AND cpu_0_instruction_master_read;
  --cpu_0/data_master granted cpu_0/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpu_0_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module))))));
    end if;

  end process;

  --cpu_0_data_master_continuerequest continued request, which is an e_mux
  cpu_0_data_master_continuerequest <= last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module AND internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  internal_cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module <= internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module AND NOT (cpu_0_data_master_arbiterlock);
  --allow new arb cycle for cpu_0/jtag_debug_module, which is an e_assign
  cpu_0_jtag_debug_module_allow_new_arb_cycle <= NOT cpu_0_data_master_arbiterlock AND NOT cpu_0_instruction_master_arbiterlock;
  --cpu_0/instruction_master assignment into master qualified-requests vector for cpu_0/jtag_debug_module, which is an e_assign
  cpu_0_jtag_debug_module_master_qreq_vector(0) <= internal_cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  --cpu_0/instruction_master grant cpu_0/jtag_debug_module, which is an e_assign
  internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module <= cpu_0_jtag_debug_module_grant_vector(0);
  --cpu_0/instruction_master saved-grant cpu_0/jtag_debug_module, which is an e_assign
  cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module <= cpu_0_jtag_debug_module_arb_winner(0) AND internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  --cpu_0/data_master assignment into master qualified-requests vector for cpu_0/jtag_debug_module, which is an e_assign
  cpu_0_jtag_debug_module_master_qreq_vector(1) <= internal_cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  --cpu_0/data_master grant cpu_0/jtag_debug_module, which is an e_assign
  internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module <= cpu_0_jtag_debug_module_grant_vector(1);
  --cpu_0/data_master saved-grant cpu_0/jtag_debug_module, which is an e_assign
  cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module <= cpu_0_jtag_debug_module_arb_winner(1) AND internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  --cpu_0/jtag_debug_module chosen-master double-vector, which is an e_assign
  cpu_0_jtag_debug_module_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((cpu_0_jtag_debug_module_master_qreq_vector & cpu_0_jtag_debug_module_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT cpu_0_jtag_debug_module_master_qreq_vector & NOT cpu_0_jtag_debug_module_master_qreq_vector))) + (std_logic_vector'("000") & (cpu_0_jtag_debug_module_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  cpu_0_jtag_debug_module_arb_winner <= A_WE_StdLogicVector((std_logic'(((cpu_0_jtag_debug_module_allow_new_arb_cycle AND or_reduce(cpu_0_jtag_debug_module_grant_vector)))) = '1'), cpu_0_jtag_debug_module_grant_vector, cpu_0_jtag_debug_module_saved_chosen_master_vector);
  --saved cpu_0_jtag_debug_module_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_jtag_debug_module_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_0_jtag_debug_module_allow_new_arb_cycle) = '1' then 
        cpu_0_jtag_debug_module_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(cpu_0_jtag_debug_module_grant_vector)) = '1'), cpu_0_jtag_debug_module_grant_vector, cpu_0_jtag_debug_module_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  cpu_0_jtag_debug_module_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((cpu_0_jtag_debug_module_chosen_master_double_vector(1) OR cpu_0_jtag_debug_module_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((cpu_0_jtag_debug_module_chosen_master_double_vector(0) OR cpu_0_jtag_debug_module_chosen_master_double_vector(2)))));
  --cpu_0/jtag_debug_module chosen master rotated left, which is an e_assign
  cpu_0_jtag_debug_module_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(cpu_0_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(cpu_0_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --cpu_0/jtag_debug_module's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_jtag_debug_module_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(cpu_0_jtag_debug_module_grant_vector)) = '1' then 
        cpu_0_jtag_debug_module_arb_addend <= A_WE_StdLogicVector((std_logic'(cpu_0_jtag_debug_module_end_xfer) = '1'), cpu_0_jtag_debug_module_chosen_master_rot_left, cpu_0_jtag_debug_module_grant_vector);
      end if;
    end if;

  end process;

  cpu_0_jtag_debug_module_begintransfer <= cpu_0_jtag_debug_module_begins_xfer;
  --cpu_0_jtag_debug_module_reset_n assignment, which is an e_assign
  cpu_0_jtag_debug_module_reset_n <= reset_n;
  --assign cpu_0_jtag_debug_module_resetrequest_from_sa = cpu_0_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_0_jtag_debug_module_resetrequest_from_sa <= cpu_0_jtag_debug_module_resetrequest;
  cpu_0_jtag_debug_module_chipselect <= internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module OR internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  --cpu_0_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  cpu_0_jtag_debug_module_firsttransfer <= A_WE_StdLogic((std_logic'(cpu_0_jtag_debug_module_begins_xfer) = '1'), cpu_0_jtag_debug_module_unreg_firsttransfer, cpu_0_jtag_debug_module_reg_firsttransfer);
  --cpu_0_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  cpu_0_jtag_debug_module_unreg_firsttransfer <= NOT ((cpu_0_jtag_debug_module_slavearbiterlockenable AND cpu_0_jtag_debug_module_any_continuerequest));
  --cpu_0_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_jtag_debug_module_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_0_jtag_debug_module_begins_xfer) = '1' then 
        cpu_0_jtag_debug_module_reg_firsttransfer <= cpu_0_jtag_debug_module_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cpu_0_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cpu_0_jtag_debug_module_beginbursttransfer_internal <= cpu_0_jtag_debug_module_begins_xfer;
  --cpu_0_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  cpu_0_jtag_debug_module_arbitration_holdoff_internal <= cpu_0_jtag_debug_module_begins_xfer AND cpu_0_jtag_debug_module_firsttransfer;
  --cpu_0_jtag_debug_module_write assignment, which is an e_mux
  cpu_0_jtag_debug_module_write <= internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module AND cpu_0_data_master_write;
  shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --cpu_0_jtag_debug_module_address mux, which is an e_mux
  cpu_0_jtag_debug_module_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module)) = '1'), (A_SRL(shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 9);
  shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master <= cpu_0_instruction_master_address_to_slave;
  --d1_cpu_0_jtag_debug_module_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cpu_0_jtag_debug_module_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cpu_0_jtag_debug_module_end_xfer <= cpu_0_jtag_debug_module_end_xfer;
    end if;

  end process;

  --cpu_0_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  cpu_0_jtag_debug_module_waits_for_read <= cpu_0_jtag_debug_module_in_a_read_cycle AND cpu_0_jtag_debug_module_begins_xfer;
  --cpu_0_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  cpu_0_jtag_debug_module_in_a_read_cycle <= ((internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module AND cpu_0_data_master_read)) OR ((internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module AND cpu_0_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cpu_0_jtag_debug_module_in_a_read_cycle;
  --cpu_0_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  cpu_0_jtag_debug_module_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_jtag_debug_module_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --cpu_0_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  cpu_0_jtag_debug_module_in_a_write_cycle <= internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cpu_0_jtag_debug_module_in_a_write_cycle;
  wait_for_cpu_0_jtag_debug_module_counter <= std_logic'('0');
  --cpu_0_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  cpu_0_jtag_debug_module_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --debugaccess mux, which is an e_mux
  cpu_0_jtag_debug_module_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_cpu_0_jtag_debug_module <= internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module <= internal_cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_cpu_0_jtag_debug_module <= internal_cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_granted_cpu_0_jtag_debug_module <= internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module <= internal_cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_requests_cpu_0_jtag_debug_module <= internal_cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
--synthesis translate_off
    --cpu_0/jtag_debug_module enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line7 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_data_master_granted_cpu_0_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_instruction_master_granted_cpu_0_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line7, now);
          write(write_line7, string'(": "));
          write(write_line7, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line7.all);
          deallocate (write_line7);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line8 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line8, now);
          write(write_line8, string'(": "));
          write(write_line8, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line8.all);
          deallocate (write_line8);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity high_res_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity high_res_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module;


architecture europa of high_res_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module;


architecture europa of jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sys_clk_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity sys_clk_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module;


architecture europa of sys_clk_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cpu_0_data_master_arbitrator is 
        port (
              -- inputs:
                 signal ad7928_spi_control_port_irq_from_sa : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_0_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal cpu_0_data_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_data_master_granted_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_gpib_edm1_clock_0_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_gpib_edm1_clock_1_in : IN STD_LOGIC;
                 signal cpu_0_data_master_granted_onchip_memory_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in : IN STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_onchip_memory_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_gpib_edm1_clock_0_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_gpib_edm1_clock_1_in : IN STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_onchip_memory_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_gpib_edm1_clock_0_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_gpib_edm1_clock_1_in : IN STD_LOGIC;
                 signal cpu_0_data_master_requests_onchip_memory_s1 : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_clk : IN STD_LOGIC;
                 signal cpu_clk_reset_n : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal d1_clock_crossing_0_s1_end_xfer : IN STD_LOGIC;
                 signal d1_cpu_0_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_cpu_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal d1_flash_ssram_pipeline_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal d1_gpib_edm1_clock_0_in_end_xfer : IN STD_LOGIC;
                 signal d1_gpib_edm1_clock_1_in_end_xfer : IN STD_LOGIC;
                 signal d1_onchip_memory_s1_end_xfer : IN STD_LOGIC;
                 signal dac_ad5308_spi_control_port_irq_from_sa : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpib_edm1_clock_1_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal high_res_timer_s1_irq_from_sa : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                 signal onchip_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal registered_cpu_0_data_master_read_data_valid_onchip_memory_s1 : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_s1_irq_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_data_master_waitrequest : OUT STD_LOGIC
              );
end entity cpu_0_data_master_arbitrator;


architecture europa of cpu_0_data_master_arbitrator is
component high_res_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component high_res_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module;

component jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module;

component sys_clk_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component sys_clk_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module;

                signal cpu_0_data_master_run :  STD_LOGIC;
                signal cpu_clk_high_res_timer_s1_irq_from_sa :  STD_LOGIC;
                signal cpu_clk_jtag_uart_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal cpu_clk_sys_clk_s1_irq_from_sa :  STD_LOGIC;
                signal internal_cpu_0_data_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal internal_cpu_0_data_master_waitrequest :  STD_LOGIC;
                signal p1_registered_cpu_0_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal registered_cpu_0_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_0_data_master_qualified_request_clock_crossing_0_s1 OR cpu_0_data_master_read_data_valid_clock_crossing_0_s1) OR NOT cpu_0_data_master_requests_clock_crossing_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_granted_clock_crossing_0_s1 OR NOT cpu_0_data_master_qualified_request_clock_crossing_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_0_data_master_qualified_request_clock_crossing_0_s1 OR NOT cpu_0_data_master_read) OR ((cpu_0_data_master_read_data_valid_clock_crossing_0_s1 AND cpu_0_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_clock_crossing_0_s1 OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT clock_crossing_0_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module OR NOT cpu_0_data_master_requests_cpu_0_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_granted_cpu_0_jtag_debug_module OR NOT cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module OR NOT cpu_0_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module OR NOT cpu_0_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 OR cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1) OR NOT cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 OR NOT cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 OR NOT cpu_0_data_master_read) OR ((cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 AND cpu_0_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT cpu_ddr_clock_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 OR cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1) OR NOT cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 OR NOT cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 OR NOT cpu_0_data_master_read) OR ((cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1 AND cpu_0_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT flash_ssram_pipeline_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_0_data_master_run <= (r_0 AND r_1) AND r_2;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in OR NOT cpu_0_data_master_requests_gpib_edm1_clock_0_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT gpib_edm1_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT gpib_edm1_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in OR NOT cpu_0_data_master_requests_gpib_edm1_clock_1_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT gpib_edm1_clock_1_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT gpib_edm1_clock_1_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_0_data_master_qualified_request_onchip_memory_s1 OR registered_cpu_0_data_master_read_data_valid_onchip_memory_s1) OR NOT cpu_0_data_master_requests_onchip_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_granted_onchip_memory_s1 OR NOT cpu_0_data_master_qualified_request_onchip_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_0_data_master_qualified_request_onchip_memory_s1 OR NOT cpu_0_data_master_read) OR ((registered_cpu_0_data_master_read_data_valid_onchip_memory_s1 AND cpu_0_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_data_master_qualified_request_onchip_memory_s1 OR NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_read OR cpu_0_data_master_write)))))))))));
  --irq assign, which is an e_assign
  cpu_0_data_master_irq <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(dac_ad5308_spi_control_port_irq_from_sa) & A_ToStdLogicVector(ad7928_spi_control_port_irq_from_sa) & A_ToStdLogicVector(cpu_clk_high_res_timer_s1_irq_from_sa) & A_ToStdLogicVector(cpu_clk_sys_clk_s1_irq_from_sa) & A_ToStdLogicVector(cpu_clk_jtag_uart_avalon_jtag_slave_irq_from_sa));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_0_data_master_address_to_slave <= cpu_0_data_master_address(27 DOWNTO 0);
  --unpredictable registered wait state incoming data, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      registered_cpu_0_data_master_readdata <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      registered_cpu_0_data_master_readdata <= p1_registered_cpu_0_data_master_readdata;
    end if;

  end process;

  --registered readdata mux, which is an e_mux
  p1_registered_cpu_0_data_master_readdata <= (((((A_REP(NOT cpu_0_data_master_requests_clock_crossing_0_s1, 32) OR clock_crossing_0_s1_readdata_from_sa)) AND ((A_REP(NOT cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1, 32) OR cpu_ddr_clock_bridge_s1_readdata_from_sa))) AND ((A_REP(NOT cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1, 32) OR flash_ssram_pipeline_bridge_s1_readdata_from_sa))) AND ((A_REP(NOT cpu_0_data_master_requests_gpib_edm1_clock_0_in, 32) OR (std_logic_vector'("0000000000000000") & (gpib_edm1_clock_0_in_readdata_from_sa))))) AND ((A_REP(NOT cpu_0_data_master_requests_gpib_edm1_clock_1_in, 32) OR gpib_edm1_clock_1_in_readdata_from_sa));
  --cpu_0/data_master readdata mux, which is an e_mux
  cpu_0_data_master_readdata <= (((((((A_REP(NOT cpu_0_data_master_requests_clock_crossing_0_s1, 32) OR registered_cpu_0_data_master_readdata)) AND ((A_REP(NOT cpu_0_data_master_requests_cpu_0_jtag_debug_module, 32) OR cpu_0_jtag_debug_module_readdata_from_sa))) AND ((A_REP(NOT cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1, 32) OR registered_cpu_0_data_master_readdata))) AND ((A_REP(NOT cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1, 32) OR registered_cpu_0_data_master_readdata))) AND ((A_REP(NOT cpu_0_data_master_requests_gpib_edm1_clock_0_in, 32) OR registered_cpu_0_data_master_readdata))) AND ((A_REP(NOT cpu_0_data_master_requests_gpib_edm1_clock_1_in, 32) OR registered_cpu_0_data_master_readdata))) AND ((A_REP(NOT cpu_0_data_master_requests_onchip_memory_s1, 32) OR onchip_memory_s1_readdata_from_sa));
  --actual waitrequest port, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_0_data_master_waitrequest <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      internal_cpu_0_data_master_waitrequest <= Vector_To_Std_Logic(NOT (A_WE_StdLogicVector((std_logic'((NOT ((cpu_0_data_master_read OR cpu_0_data_master_write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_data_master_run AND internal_cpu_0_data_master_waitrequest))))))));
    end if;

  end process;

  --high_res_timer_s1_irq_from_sa from pll_c2_out to cpu_clk
  high_res_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master : high_res_timer_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module
    port map(
      data_out => cpu_clk_high_res_timer_s1_irq_from_sa,
      clk => cpu_clk,
      data_in => high_res_timer_s1_irq_from_sa,
      reset_n => cpu_clk_reset_n
    );


  --jtag_uart_avalon_jtag_slave_irq_from_sa from pll_c2_out to cpu_clk
  jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master : jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_0_data_master_module
    port map(
      data_out => cpu_clk_jtag_uart_avalon_jtag_slave_irq_from_sa,
      clk => cpu_clk,
      data_in => jtag_uart_avalon_jtag_slave_irq_from_sa,
      reset_n => cpu_clk_reset_n
    );


  --sys_clk_s1_irq_from_sa from pll_c2_out to cpu_clk
  sys_clk_s1_irq_from_sa_clock_crossing_cpu_0_data_master : sys_clk_s1_irq_from_sa_clock_crossing_cpu_0_data_master_module
    port map(
      data_out => cpu_clk_sys_clk_s1_irq_from_sa,
      clk => cpu_clk,
      data_in => sys_clk_s1_irq_from_sa,
      reset_n => cpu_clk_reset_n
    );


  --vhdl renameroo for output signals
  cpu_0_data_master_address_to_slave <= internal_cpu_0_data_master_address_to_slave;
  --vhdl renameroo for output signals
  cpu_0_data_master_waitrequest <= internal_cpu_0_data_master_waitrequest;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_0_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_0_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal cpu_0_instruction_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_instruction_master_granted_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_granted_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_granted_onchip_memory_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_onchip_memory_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_onchip_memory_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_requests_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_requests_cpu_0_jtag_debug_module : IN STD_LOGIC;
                 signal cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_0_instruction_master_requests_onchip_memory_s1 : IN STD_LOGIC;
                 signal cpu_0_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal d1_clock_crossing_0_s1_end_xfer : IN STD_LOGIC;
                 signal d1_cpu_0_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_cpu_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal d1_flash_ssram_pipeline_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal d1_onchip_memory_s1_end_xfer : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal onchip_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_instruction_master_waitrequest : OUT STD_LOGIC
              );
end entity cpu_0_instruction_master_arbitrator;


architecture europa of cpu_0_instruction_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpu_0_instruction_master_address_last_time :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_0_instruction_master_read_last_time :  STD_LOGIC;
                signal cpu_0_instruction_master_run :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal internal_cpu_0_instruction_master_waitrequest :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 OR cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1) OR NOT cpu_0_instruction_master_requests_clock_crossing_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_instruction_master_granted_clock_crossing_0_s1 OR NOT cpu_0_instruction_master_qualified_request_clock_crossing_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 OR NOT cpu_0_instruction_master_read) OR ((cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1 AND cpu_0_instruction_master_read)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module OR NOT cpu_0_instruction_master_requests_cpu_0_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_instruction_master_granted_cpu_0_jtag_debug_module OR NOT cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module OR NOT cpu_0_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cpu_0_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_read)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 OR cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1) OR NOT cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 OR NOT cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 OR NOT cpu_0_instruction_master_read) OR ((cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 AND cpu_0_instruction_master_read)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 OR cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1) OR NOT cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 OR NOT cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 OR NOT cpu_0_instruction_master_read) OR ((cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1 AND cpu_0_instruction_master_read)))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_0_instruction_master_run <= r_0 AND r_2;
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpu_0_instruction_master_qualified_request_onchip_memory_s1 OR cpu_0_instruction_master_read_data_valid_onchip_memory_s1) OR NOT cpu_0_instruction_master_requests_onchip_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_0_instruction_master_granted_onchip_memory_s1 OR NOT cpu_0_instruction_master_qualified_request_onchip_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpu_0_instruction_master_qualified_request_onchip_memory_s1 OR NOT cpu_0_instruction_master_read) OR ((cpu_0_instruction_master_read_data_valid_onchip_memory_s1 AND cpu_0_instruction_master_read)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_0_instruction_master_address_to_slave <= cpu_0_instruction_master_address(27 DOWNTO 0);
  --cpu_0/instruction_master readdata mux, which is an e_mux
  cpu_0_instruction_master_readdata <= (((((A_REP(NOT cpu_0_instruction_master_requests_clock_crossing_0_s1, 32) OR clock_crossing_0_s1_readdata_from_sa)) AND ((A_REP(NOT cpu_0_instruction_master_requests_cpu_0_jtag_debug_module, 32) OR cpu_0_jtag_debug_module_readdata_from_sa))) AND ((A_REP(NOT cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1, 32) OR cpu_ddr_clock_bridge_s1_readdata_from_sa))) AND ((A_REP(NOT cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1, 32) OR flash_ssram_pipeline_bridge_s1_readdata_from_sa))) AND ((A_REP(NOT cpu_0_instruction_master_requests_onchip_memory_s1, 32) OR onchip_memory_s1_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_cpu_0_instruction_master_waitrequest <= NOT cpu_0_instruction_master_run;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_address_to_slave <= internal_cpu_0_instruction_master_address_to_slave;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_waitrequest <= internal_cpu_0_instruction_master_waitrequest;
--synthesis translate_off
    --cpu_0_instruction_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_0_instruction_master_address_last_time <= std_logic_vector'("0000000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_0_instruction_master_address_last_time <= cpu_0_instruction_master_address;
      end if;

    end process;

    --cpu_0/instruction_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpu_0_instruction_master_waitrequest AND (cpu_0_instruction_master_read);
      end if;

    end process;

    --cpu_0_instruction_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line9 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_0_instruction_master_address /= cpu_0_instruction_master_address_last_time))))) = '1' then 
          write(write_line9, now);
          write(write_line9, string'(": "));
          write(write_line9, string'("cpu_0_instruction_master_address did not heed wait!!!"));
          write(output, write_line9.all);
          deallocate (write_line9);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_0_instruction_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_0_instruction_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_0_instruction_master_read_last_time <= cpu_0_instruction_master_read;
      end if;

    end process;

    --cpu_0_instruction_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line10 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_0_instruction_master_read) /= std_logic'(cpu_0_instruction_master_read_last_time)))))) = '1' then 
          write(write_line10, now);
          write(write_line10, string'(": "));
          write(write_line10, string'("cpu_0_instruction_master_read did not heed wait!!!"));
          write(output, write_line10.all);
          deallocate (write_line10);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_0_data_master_to_cpu_ddr_clock_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_0_data_master_to_cpu_ddr_clock_bridge_s1_module;


architecture europa of rdv_fifo_for_cpu_0_data_master_to_cpu_ddr_clock_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_33 :  STD_LOGIC;
                signal full_34 :  STD_LOGIC;
                signal full_35 :  STD_LOGIC;
                signal full_36 :  STD_LOGIC;
                signal full_37 :  STD_LOGIC;
                signal full_38 :  STD_LOGIC;
                signal full_39 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_40 :  STD_LOGIC;
                signal full_41 :  STD_LOGIC;
                signal full_42 :  STD_LOGIC;
                signal full_43 :  STD_LOGIC;
                signal full_44 :  STD_LOGIC;
                signal full_45 :  STD_LOGIC;
                signal full_46 :  STD_LOGIC;
                signal full_47 :  STD_LOGIC;
                signal full_48 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p32_full_32 :  STD_LOGIC;
                signal p32_stage_32 :  STD_LOGIC;
                signal p33_full_33 :  STD_LOGIC;
                signal p33_stage_33 :  STD_LOGIC;
                signal p34_full_34 :  STD_LOGIC;
                signal p34_stage_34 :  STD_LOGIC;
                signal p35_full_35 :  STD_LOGIC;
                signal p35_stage_35 :  STD_LOGIC;
                signal p36_full_36 :  STD_LOGIC;
                signal p36_stage_36 :  STD_LOGIC;
                signal p37_full_37 :  STD_LOGIC;
                signal p37_stage_37 :  STD_LOGIC;
                signal p38_full_38 :  STD_LOGIC;
                signal p38_stage_38 :  STD_LOGIC;
                signal p39_full_39 :  STD_LOGIC;
                signal p39_stage_39 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p40_full_40 :  STD_LOGIC;
                signal p40_stage_40 :  STD_LOGIC;
                signal p41_full_41 :  STD_LOGIC;
                signal p41_stage_41 :  STD_LOGIC;
                signal p42_full_42 :  STD_LOGIC;
                signal p42_stage_42 :  STD_LOGIC;
                signal p43_full_43 :  STD_LOGIC;
                signal p43_stage_43 :  STD_LOGIC;
                signal p44_full_44 :  STD_LOGIC;
                signal p44_stage_44 :  STD_LOGIC;
                signal p45_full_45 :  STD_LOGIC;
                signal p45_stage_45 :  STD_LOGIC;
                signal p46_full_46 :  STD_LOGIC;
                signal p46_stage_46 :  STD_LOGIC;
                signal p47_full_47 :  STD_LOGIC;
                signal p47_stage_47 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_32 :  STD_LOGIC;
                signal stage_33 :  STD_LOGIC;
                signal stage_34 :  STD_LOGIC;
                signal stage_35 :  STD_LOGIC;
                signal stage_36 :  STD_LOGIC;
                signal stage_37 :  STD_LOGIC;
                signal stage_38 :  STD_LOGIC;
                signal stage_39 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_40 :  STD_LOGIC;
                signal stage_41 :  STD_LOGIC;
                signal stage_42 :  STD_LOGIC;
                signal stage_43 :  STD_LOGIC;
                signal stage_44 :  STD_LOGIC;
                signal stage_45 :  STD_LOGIC;
                signal stage_46 :  STD_LOGIC;
                signal stage_47 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_47;
  empty <= NOT(full_0);
  full_48 <= std_logic'('0');
  --data_47, which is an e_mux
  p47_stage_47 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_48 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_47, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_47 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_47))))) = '1' then 
        if std_logic'(((sync_reset AND full_47) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_48))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_47 <= std_logic'('0');
        else
          stage_47 <= p47_stage_47;
        end if;
      end if;
    end if;

  end process;

  --control_47, which is an e_mux
  p47_full_47 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_46))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_47, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_47 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_47 <= std_logic'('0');
        else
          full_47 <= p47_full_47;
        end if;
      end if;
    end if;

  end process;

  --data_46, which is an e_mux
  p46_stage_46 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_47 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_47);
  --data_reg_46, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_46 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_46))))) = '1' then 
        if std_logic'(((sync_reset AND full_46) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_47))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_46 <= std_logic'('0');
        else
          stage_46 <= p46_stage_46;
        end if;
      end if;
    end if;

  end process;

  --control_46, which is an e_mux
  p46_full_46 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_45, full_47);
  --control_reg_46, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_46 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_46 <= std_logic'('0');
        else
          full_46 <= p46_full_46;
        end if;
      end if;
    end if;

  end process;

  --data_45, which is an e_mux
  p45_stage_45 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_46 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_46);
  --data_reg_45, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_45 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_45))))) = '1' then 
        if std_logic'(((sync_reset AND full_45) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_46))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_45 <= std_logic'('0');
        else
          stage_45 <= p45_stage_45;
        end if;
      end if;
    end if;

  end process;

  --control_45, which is an e_mux
  p45_full_45 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_44, full_46);
  --control_reg_45, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_45 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_45 <= std_logic'('0');
        else
          full_45 <= p45_full_45;
        end if;
      end if;
    end if;

  end process;

  --data_44, which is an e_mux
  p44_stage_44 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_45 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_45);
  --data_reg_44, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_44 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_44))))) = '1' then 
        if std_logic'(((sync_reset AND full_44) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_45))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_44 <= std_logic'('0');
        else
          stage_44 <= p44_stage_44;
        end if;
      end if;
    end if;

  end process;

  --control_44, which is an e_mux
  p44_full_44 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_43, full_45);
  --control_reg_44, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_44 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_44 <= std_logic'('0');
        else
          full_44 <= p44_full_44;
        end if;
      end if;
    end if;

  end process;

  --data_43, which is an e_mux
  p43_stage_43 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_44 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_44);
  --data_reg_43, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_43 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_43))))) = '1' then 
        if std_logic'(((sync_reset AND full_43) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_44))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_43 <= std_logic'('0');
        else
          stage_43 <= p43_stage_43;
        end if;
      end if;
    end if;

  end process;

  --control_43, which is an e_mux
  p43_full_43 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_42, full_44);
  --control_reg_43, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_43 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_43 <= std_logic'('0');
        else
          full_43 <= p43_full_43;
        end if;
      end if;
    end if;

  end process;

  --data_42, which is an e_mux
  p42_stage_42 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_43 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_43);
  --data_reg_42, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_42 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_42))))) = '1' then 
        if std_logic'(((sync_reset AND full_42) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_43))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_42 <= std_logic'('0');
        else
          stage_42 <= p42_stage_42;
        end if;
      end if;
    end if;

  end process;

  --control_42, which is an e_mux
  p42_full_42 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_41, full_43);
  --control_reg_42, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_42 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_42 <= std_logic'('0');
        else
          full_42 <= p42_full_42;
        end if;
      end if;
    end if;

  end process;

  --data_41, which is an e_mux
  p41_stage_41 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_42 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_42);
  --data_reg_41, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_41 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_41))))) = '1' then 
        if std_logic'(((sync_reset AND full_41) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_42))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_41 <= std_logic'('0');
        else
          stage_41 <= p41_stage_41;
        end if;
      end if;
    end if;

  end process;

  --control_41, which is an e_mux
  p41_full_41 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_40, full_42);
  --control_reg_41, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_41 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_41 <= std_logic'('0');
        else
          full_41 <= p41_full_41;
        end if;
      end if;
    end if;

  end process;

  --data_40, which is an e_mux
  p40_stage_40 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_41 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_41);
  --data_reg_40, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_40 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_40))))) = '1' then 
        if std_logic'(((sync_reset AND full_40) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_41))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_40 <= std_logic'('0');
        else
          stage_40 <= p40_stage_40;
        end if;
      end if;
    end if;

  end process;

  --control_40, which is an e_mux
  p40_full_40 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_39, full_41);
  --control_reg_40, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_40 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_40 <= std_logic'('0');
        else
          full_40 <= p40_full_40;
        end if;
      end if;
    end if;

  end process;

  --data_39, which is an e_mux
  p39_stage_39 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_40 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_40);
  --data_reg_39, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_39 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_39))))) = '1' then 
        if std_logic'(((sync_reset AND full_39) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_40))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_39 <= std_logic'('0');
        else
          stage_39 <= p39_stage_39;
        end if;
      end if;
    end if;

  end process;

  --control_39, which is an e_mux
  p39_full_39 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_38, full_40);
  --control_reg_39, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_39 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_39 <= std_logic'('0');
        else
          full_39 <= p39_full_39;
        end if;
      end if;
    end if;

  end process;

  --data_38, which is an e_mux
  p38_stage_38 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_39 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_39);
  --data_reg_38, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_38 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_38))))) = '1' then 
        if std_logic'(((sync_reset AND full_38) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_39))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_38 <= std_logic'('0');
        else
          stage_38 <= p38_stage_38;
        end if;
      end if;
    end if;

  end process;

  --control_38, which is an e_mux
  p38_full_38 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_37, full_39);
  --control_reg_38, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_38 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_38 <= std_logic'('0');
        else
          full_38 <= p38_full_38;
        end if;
      end if;
    end if;

  end process;

  --data_37, which is an e_mux
  p37_stage_37 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_38 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_38);
  --data_reg_37, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_37 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_37))))) = '1' then 
        if std_logic'(((sync_reset AND full_37) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_38))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_37 <= std_logic'('0');
        else
          stage_37 <= p37_stage_37;
        end if;
      end if;
    end if;

  end process;

  --control_37, which is an e_mux
  p37_full_37 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_36, full_38);
  --control_reg_37, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_37 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_37 <= std_logic'('0');
        else
          full_37 <= p37_full_37;
        end if;
      end if;
    end if;

  end process;

  --data_36, which is an e_mux
  p36_stage_36 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_37 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_37);
  --data_reg_36, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_36 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_36))))) = '1' then 
        if std_logic'(((sync_reset AND full_36) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_37))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_36 <= std_logic'('0');
        else
          stage_36 <= p36_stage_36;
        end if;
      end if;
    end if;

  end process;

  --control_36, which is an e_mux
  p36_full_36 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_35, full_37);
  --control_reg_36, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_36 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_36 <= std_logic'('0');
        else
          full_36 <= p36_full_36;
        end if;
      end if;
    end if;

  end process;

  --data_35, which is an e_mux
  p35_stage_35 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_36 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_36);
  --data_reg_35, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_35 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_35))))) = '1' then 
        if std_logic'(((sync_reset AND full_35) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_36))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_35 <= std_logic'('0');
        else
          stage_35 <= p35_stage_35;
        end if;
      end if;
    end if;

  end process;

  --control_35, which is an e_mux
  p35_full_35 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_34, full_36);
  --control_reg_35, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_35 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_35 <= std_logic'('0');
        else
          full_35 <= p35_full_35;
        end if;
      end if;
    end if;

  end process;

  --data_34, which is an e_mux
  p34_stage_34 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_35 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_35);
  --data_reg_34, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_34 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_34))))) = '1' then 
        if std_logic'(((sync_reset AND full_34) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_35))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_34 <= std_logic'('0');
        else
          stage_34 <= p34_stage_34;
        end if;
      end if;
    end if;

  end process;

  --control_34, which is an e_mux
  p34_full_34 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_33, full_35);
  --control_reg_34, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_34 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_34 <= std_logic'('0');
        else
          full_34 <= p34_full_34;
        end if;
      end if;
    end if;

  end process;

  --data_33, which is an e_mux
  p33_stage_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_34 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_34);
  --data_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_33))))) = '1' then 
        if std_logic'(((sync_reset AND full_33) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_34))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_33 <= std_logic'('0');
        else
          stage_33 <= p33_stage_33;
        end if;
      end if;
    end if;

  end process;

  --control_33, which is an e_mux
  p33_full_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_32, full_34);
  --control_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_33 <= std_logic'('0');
        else
          full_33 <= p33_full_33;
        end if;
      end if;
    end if;

  end process;

  --data_32, which is an e_mux
  p32_stage_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_33 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_33);
  --data_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_32))))) = '1' then 
        if std_logic'(((sync_reset AND full_32) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_33))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_32 <= std_logic'('0');
        else
          stage_32 <= p32_stage_32;
        end if;
      end if;
    end if;

  end process;

  --control_32, which is an e_mux
  p32_full_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_31, full_33);
  --control_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_32 <= std_logic'('0');
        else
          full_32 <= p32_full_32;
        end if;
      end if;
    end if;

  end process;

  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_32);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_30, full_32);
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_0_instruction_master_to_cpu_ddr_clock_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_0_instruction_master_to_cpu_ddr_clock_bridge_s1_module;


architecture europa of rdv_fifo_for_cpu_0_instruction_master_to_cpu_ddr_clock_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_33 :  STD_LOGIC;
                signal full_34 :  STD_LOGIC;
                signal full_35 :  STD_LOGIC;
                signal full_36 :  STD_LOGIC;
                signal full_37 :  STD_LOGIC;
                signal full_38 :  STD_LOGIC;
                signal full_39 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_40 :  STD_LOGIC;
                signal full_41 :  STD_LOGIC;
                signal full_42 :  STD_LOGIC;
                signal full_43 :  STD_LOGIC;
                signal full_44 :  STD_LOGIC;
                signal full_45 :  STD_LOGIC;
                signal full_46 :  STD_LOGIC;
                signal full_47 :  STD_LOGIC;
                signal full_48 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p32_full_32 :  STD_LOGIC;
                signal p32_stage_32 :  STD_LOGIC;
                signal p33_full_33 :  STD_LOGIC;
                signal p33_stage_33 :  STD_LOGIC;
                signal p34_full_34 :  STD_LOGIC;
                signal p34_stage_34 :  STD_LOGIC;
                signal p35_full_35 :  STD_LOGIC;
                signal p35_stage_35 :  STD_LOGIC;
                signal p36_full_36 :  STD_LOGIC;
                signal p36_stage_36 :  STD_LOGIC;
                signal p37_full_37 :  STD_LOGIC;
                signal p37_stage_37 :  STD_LOGIC;
                signal p38_full_38 :  STD_LOGIC;
                signal p38_stage_38 :  STD_LOGIC;
                signal p39_full_39 :  STD_LOGIC;
                signal p39_stage_39 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p40_full_40 :  STD_LOGIC;
                signal p40_stage_40 :  STD_LOGIC;
                signal p41_full_41 :  STD_LOGIC;
                signal p41_stage_41 :  STD_LOGIC;
                signal p42_full_42 :  STD_LOGIC;
                signal p42_stage_42 :  STD_LOGIC;
                signal p43_full_43 :  STD_LOGIC;
                signal p43_stage_43 :  STD_LOGIC;
                signal p44_full_44 :  STD_LOGIC;
                signal p44_stage_44 :  STD_LOGIC;
                signal p45_full_45 :  STD_LOGIC;
                signal p45_stage_45 :  STD_LOGIC;
                signal p46_full_46 :  STD_LOGIC;
                signal p46_stage_46 :  STD_LOGIC;
                signal p47_full_47 :  STD_LOGIC;
                signal p47_stage_47 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_32 :  STD_LOGIC;
                signal stage_33 :  STD_LOGIC;
                signal stage_34 :  STD_LOGIC;
                signal stage_35 :  STD_LOGIC;
                signal stage_36 :  STD_LOGIC;
                signal stage_37 :  STD_LOGIC;
                signal stage_38 :  STD_LOGIC;
                signal stage_39 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_40 :  STD_LOGIC;
                signal stage_41 :  STD_LOGIC;
                signal stage_42 :  STD_LOGIC;
                signal stage_43 :  STD_LOGIC;
                signal stage_44 :  STD_LOGIC;
                signal stage_45 :  STD_LOGIC;
                signal stage_46 :  STD_LOGIC;
                signal stage_47 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_47;
  empty <= NOT(full_0);
  full_48 <= std_logic'('0');
  --data_47, which is an e_mux
  p47_stage_47 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_48 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_47, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_47 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_47))))) = '1' then 
        if std_logic'(((sync_reset AND full_47) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_48))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_47 <= std_logic'('0');
        else
          stage_47 <= p47_stage_47;
        end if;
      end if;
    end if;

  end process;

  --control_47, which is an e_mux
  p47_full_47 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_46))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_47, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_47 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_47 <= std_logic'('0');
        else
          full_47 <= p47_full_47;
        end if;
      end if;
    end if;

  end process;

  --data_46, which is an e_mux
  p46_stage_46 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_47 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_47);
  --data_reg_46, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_46 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_46))))) = '1' then 
        if std_logic'(((sync_reset AND full_46) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_47))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_46 <= std_logic'('0');
        else
          stage_46 <= p46_stage_46;
        end if;
      end if;
    end if;

  end process;

  --control_46, which is an e_mux
  p46_full_46 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_45, full_47);
  --control_reg_46, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_46 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_46 <= std_logic'('0');
        else
          full_46 <= p46_full_46;
        end if;
      end if;
    end if;

  end process;

  --data_45, which is an e_mux
  p45_stage_45 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_46 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_46);
  --data_reg_45, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_45 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_45))))) = '1' then 
        if std_logic'(((sync_reset AND full_45) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_46))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_45 <= std_logic'('0');
        else
          stage_45 <= p45_stage_45;
        end if;
      end if;
    end if;

  end process;

  --control_45, which is an e_mux
  p45_full_45 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_44, full_46);
  --control_reg_45, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_45 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_45 <= std_logic'('0');
        else
          full_45 <= p45_full_45;
        end if;
      end if;
    end if;

  end process;

  --data_44, which is an e_mux
  p44_stage_44 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_45 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_45);
  --data_reg_44, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_44 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_44))))) = '1' then 
        if std_logic'(((sync_reset AND full_44) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_45))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_44 <= std_logic'('0');
        else
          stage_44 <= p44_stage_44;
        end if;
      end if;
    end if;

  end process;

  --control_44, which is an e_mux
  p44_full_44 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_43, full_45);
  --control_reg_44, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_44 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_44 <= std_logic'('0');
        else
          full_44 <= p44_full_44;
        end if;
      end if;
    end if;

  end process;

  --data_43, which is an e_mux
  p43_stage_43 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_44 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_44);
  --data_reg_43, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_43 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_43))))) = '1' then 
        if std_logic'(((sync_reset AND full_43) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_44))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_43 <= std_logic'('0');
        else
          stage_43 <= p43_stage_43;
        end if;
      end if;
    end if;

  end process;

  --control_43, which is an e_mux
  p43_full_43 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_42, full_44);
  --control_reg_43, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_43 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_43 <= std_logic'('0');
        else
          full_43 <= p43_full_43;
        end if;
      end if;
    end if;

  end process;

  --data_42, which is an e_mux
  p42_stage_42 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_43 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_43);
  --data_reg_42, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_42 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_42))))) = '1' then 
        if std_logic'(((sync_reset AND full_42) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_43))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_42 <= std_logic'('0');
        else
          stage_42 <= p42_stage_42;
        end if;
      end if;
    end if;

  end process;

  --control_42, which is an e_mux
  p42_full_42 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_41, full_43);
  --control_reg_42, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_42 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_42 <= std_logic'('0');
        else
          full_42 <= p42_full_42;
        end if;
      end if;
    end if;

  end process;

  --data_41, which is an e_mux
  p41_stage_41 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_42 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_42);
  --data_reg_41, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_41 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_41))))) = '1' then 
        if std_logic'(((sync_reset AND full_41) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_42))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_41 <= std_logic'('0');
        else
          stage_41 <= p41_stage_41;
        end if;
      end if;
    end if;

  end process;

  --control_41, which is an e_mux
  p41_full_41 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_40, full_42);
  --control_reg_41, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_41 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_41 <= std_logic'('0');
        else
          full_41 <= p41_full_41;
        end if;
      end if;
    end if;

  end process;

  --data_40, which is an e_mux
  p40_stage_40 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_41 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_41);
  --data_reg_40, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_40 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_40))))) = '1' then 
        if std_logic'(((sync_reset AND full_40) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_41))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_40 <= std_logic'('0');
        else
          stage_40 <= p40_stage_40;
        end if;
      end if;
    end if;

  end process;

  --control_40, which is an e_mux
  p40_full_40 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_39, full_41);
  --control_reg_40, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_40 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_40 <= std_logic'('0');
        else
          full_40 <= p40_full_40;
        end if;
      end if;
    end if;

  end process;

  --data_39, which is an e_mux
  p39_stage_39 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_40 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_40);
  --data_reg_39, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_39 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_39))))) = '1' then 
        if std_logic'(((sync_reset AND full_39) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_40))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_39 <= std_logic'('0');
        else
          stage_39 <= p39_stage_39;
        end if;
      end if;
    end if;

  end process;

  --control_39, which is an e_mux
  p39_full_39 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_38, full_40);
  --control_reg_39, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_39 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_39 <= std_logic'('0');
        else
          full_39 <= p39_full_39;
        end if;
      end if;
    end if;

  end process;

  --data_38, which is an e_mux
  p38_stage_38 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_39 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_39);
  --data_reg_38, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_38 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_38))))) = '1' then 
        if std_logic'(((sync_reset AND full_38) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_39))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_38 <= std_logic'('0');
        else
          stage_38 <= p38_stage_38;
        end if;
      end if;
    end if;

  end process;

  --control_38, which is an e_mux
  p38_full_38 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_37, full_39);
  --control_reg_38, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_38 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_38 <= std_logic'('0');
        else
          full_38 <= p38_full_38;
        end if;
      end if;
    end if;

  end process;

  --data_37, which is an e_mux
  p37_stage_37 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_38 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_38);
  --data_reg_37, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_37 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_37))))) = '1' then 
        if std_logic'(((sync_reset AND full_37) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_38))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_37 <= std_logic'('0');
        else
          stage_37 <= p37_stage_37;
        end if;
      end if;
    end if;

  end process;

  --control_37, which is an e_mux
  p37_full_37 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_36, full_38);
  --control_reg_37, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_37 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_37 <= std_logic'('0');
        else
          full_37 <= p37_full_37;
        end if;
      end if;
    end if;

  end process;

  --data_36, which is an e_mux
  p36_stage_36 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_37 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_37);
  --data_reg_36, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_36 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_36))))) = '1' then 
        if std_logic'(((sync_reset AND full_36) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_37))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_36 <= std_logic'('0');
        else
          stage_36 <= p36_stage_36;
        end if;
      end if;
    end if;

  end process;

  --control_36, which is an e_mux
  p36_full_36 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_35, full_37);
  --control_reg_36, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_36 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_36 <= std_logic'('0');
        else
          full_36 <= p36_full_36;
        end if;
      end if;
    end if;

  end process;

  --data_35, which is an e_mux
  p35_stage_35 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_36 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_36);
  --data_reg_35, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_35 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_35))))) = '1' then 
        if std_logic'(((sync_reset AND full_35) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_36))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_35 <= std_logic'('0');
        else
          stage_35 <= p35_stage_35;
        end if;
      end if;
    end if;

  end process;

  --control_35, which is an e_mux
  p35_full_35 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_34, full_36);
  --control_reg_35, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_35 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_35 <= std_logic'('0');
        else
          full_35 <= p35_full_35;
        end if;
      end if;
    end if;

  end process;

  --data_34, which is an e_mux
  p34_stage_34 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_35 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_35);
  --data_reg_34, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_34 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_34))))) = '1' then 
        if std_logic'(((sync_reset AND full_34) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_35))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_34 <= std_logic'('0');
        else
          stage_34 <= p34_stage_34;
        end if;
      end if;
    end if;

  end process;

  --control_34, which is an e_mux
  p34_full_34 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_33, full_35);
  --control_reg_34, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_34 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_34 <= std_logic'('0');
        else
          full_34 <= p34_full_34;
        end if;
      end if;
    end if;

  end process;

  --data_33, which is an e_mux
  p33_stage_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_34 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_34);
  --data_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_33))))) = '1' then 
        if std_logic'(((sync_reset AND full_33) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_34))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_33 <= std_logic'('0');
        else
          stage_33 <= p33_stage_33;
        end if;
      end if;
    end if;

  end process;

  --control_33, which is an e_mux
  p33_full_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_32, full_34);
  --control_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_33 <= std_logic'('0');
        else
          full_33 <= p33_full_33;
        end if;
      end if;
    end if;

  end process;

  --data_32, which is an e_mux
  p32_stage_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_33 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_33);
  --data_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_32))))) = '1' then 
        if std_logic'(((sync_reset AND full_32) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_33))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_32 <= std_logic'('0');
        else
          stage_32 <= p32_stage_32;
        end if;
      end if;
    end if;

  end process;

  --control_32, which is an e_mux
  p32_full_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_31, full_33);
  --control_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_32 <= std_logic'('0');
        else
          full_32 <= p32_full_32;
        end if;
      end if;
    end if;

  end process;

  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_32);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_30, full_32);
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_ddr_clock_bridge_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_instruction_master_read : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_endofpacket : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_readdatavalid : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_read : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_reset_n : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_write : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_ddr_clock_bridge_s1_end_xfer : OUT STD_LOGIC
              );
end entity cpu_ddr_clock_bridge_s1_arbitrator;


architecture europa of cpu_ddr_clock_bridge_s1_arbitrator is
component rdv_fifo_for_cpu_0_data_master_to_cpu_ddr_clock_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_0_data_master_to_cpu_ddr_clock_bridge_s1_module;

component rdv_fifo_for_cpu_0_instruction_master_to_cpu_ddr_clock_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_0_instruction_master_to_cpu_ddr_clock_bridge_s1_module;

                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_0_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_allgrants :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_any_continuerequest :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_arb_counter_enable :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_arb_share_counter :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_arb_share_set_values :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_begins_xfer :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_end_xfer :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_firsttransfer :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_in_a_read_cycle :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_in_a_write_cycle :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_non_bursting_master_requests :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_reg_firsttransfer :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_slavearbiterlockenable :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_unreg_firsttransfer :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_waits_for_read :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_cpu_0_data_master_granted_slave_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal last_cycle_cpu_0_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal module_input10 :  STD_LOGIC;
                signal module_input11 :  STD_LOGIC;
                signal module_input6 :  STD_LOGIC;
                signal module_input7 :  STD_LOGIC;
                signal module_input8 :  STD_LOGIC;
                signal module_input9 :  STD_LOGIC;
                signal shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_0_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_0_instruction_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_cpu_ddr_clock_bridge_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cpu_ddr_clock_bridge_s1_end_xfer;
    end if;

  end process;

  cpu_ddr_clock_bridge_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 OR internal_cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1));
  --assign cpu_ddr_clock_bridge_s1_readdata_from_sa = cpu_ddr_clock_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_ddr_clock_bridge_s1_readdata_from_sa <= cpu_ddr_clock_bridge_s1_readdata;
  internal_cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(27 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("0100000000000000000000000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign cpu_ddr_clock_bridge_s1_waitrequest_from_sa = cpu_ddr_clock_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_cpu_ddr_clock_bridge_s1_waitrequest_from_sa <= cpu_ddr_clock_bridge_s1_waitrequest;
  --assign cpu_ddr_clock_bridge_s1_readdatavalid_from_sa = cpu_ddr_clock_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_ddr_clock_bridge_s1_readdatavalid_from_sa <= cpu_ddr_clock_bridge_s1_readdatavalid;
  --cpu_ddr_clock_bridge_s1_arb_share_counter set values, which is an e_mux
  cpu_ddr_clock_bridge_s1_arb_share_set_values <= std_logic'('1');
  --cpu_ddr_clock_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_non_bursting_master_requests <= ((internal_cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 OR internal_cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1) OR internal_cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1) OR internal_cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  --cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --cpu_ddr_clock_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  cpu_ddr_clock_bridge_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_ddr_clock_bridge_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(cpu_ddr_clock_bridge_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --cpu_ddr_clock_bridge_s1_allgrants all slave grants, which is an e_mux
  cpu_ddr_clock_bridge_s1_allgrants <= (((or_reduce(cpu_ddr_clock_bridge_s1_grant_vector)) OR (or_reduce(cpu_ddr_clock_bridge_s1_grant_vector))) OR (or_reduce(cpu_ddr_clock_bridge_s1_grant_vector))) OR (or_reduce(cpu_ddr_clock_bridge_s1_grant_vector));
  --cpu_ddr_clock_bridge_s1_end_xfer assignment, which is an e_assign
  cpu_ddr_clock_bridge_s1_end_xfer <= NOT ((cpu_ddr_clock_bridge_s1_waits_for_read OR cpu_ddr_clock_bridge_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 <= cpu_ddr_clock_bridge_s1_end_xfer AND (((NOT cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cpu_ddr_clock_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  cpu_ddr_clock_bridge_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 AND cpu_ddr_clock_bridge_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 AND NOT cpu_ddr_clock_bridge_s1_non_bursting_master_requests));
  --cpu_ddr_clock_bridge_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_ddr_clock_bridge_s1_arb_counter_enable) = '1' then 
        cpu_ddr_clock_bridge_s1_arb_share_counter <= cpu_ddr_clock_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_ddr_clock_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(cpu_ddr_clock_bridge_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1)) OR ((end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 AND NOT cpu_ddr_clock_bridge_s1_non_bursting_master_requests)))) = '1' then 
        cpu_ddr_clock_bridge_s1_slavearbiterlockenable <= cpu_ddr_clock_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_0/data_master cpu_ddr_clock_bridge/s1 arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= cpu_ddr_clock_bridge_s1_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 <= cpu_ddr_clock_bridge_s1_arb_share_counter_next_value;
  --cpu_0/data_master cpu_ddr_clock_bridge/s1 arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --cpu_0/instruction_master cpu_ddr_clock_bridge/s1 arbiterlock, which is an e_assign
  cpu_0_instruction_master_arbiterlock <= cpu_ddr_clock_bridge_s1_slavearbiterlockenable AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master cpu_ddr_clock_bridge/s1 arbiterlock2, which is an e_assign
  cpu_0_instruction_master_arbiterlock2 <= cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master granted cpu_ddr_clock_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal OR NOT internal_cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1))))));
    end if;

  end process;

  --cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  cpu_0_instruction_master_continuerequest <= last_cycle_cpu_0_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 AND internal_cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  --cpu_ddr_clock_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  cpu_ddr_clock_bridge_s1_any_continuerequest <= cpu_0_instruction_master_continuerequest OR cpu_0_data_master_continuerequest;
  internal_cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 <= internal_cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 AND NOT (((((cpu_0_data_master_read AND ((NOT cpu_0_data_master_waitrequest OR (internal_cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register))))) OR (((NOT cpu_0_data_master_waitrequest) AND cpu_0_data_master_write))) OR cpu_0_instruction_master_arbiterlock));
  --unique name for cpu_ddr_clock_bridge_s1_move_on_to_next_transaction, which is an e_assign
  cpu_ddr_clock_bridge_s1_move_on_to_next_transaction <= cpu_ddr_clock_bridge_s1_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_0_data_master_to_cpu_ddr_clock_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_0_data_master_to_cpu_ddr_clock_bridge_s1 : rdv_fifo_for_cpu_0_data_master_to_cpu_ddr_clock_bridge_s1_module
    port map(
      data_out => cpu_0_data_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1,
      empty => open,
      fifo_contains_ones_n => cpu_0_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1,
      full => open,
      clear_fifo => module_input6,
      clk => clk,
      data_in => internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1,
      read => cpu_ddr_clock_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input7,
      write => module_input8
    );

  module_input6 <= std_logic'('0');
  module_input7 <= std_logic'('0');
  module_input8 <= in_a_read_cycle AND NOT cpu_ddr_clock_bridge_s1_waits_for_read;

  internal_cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register <= NOT cpu_0_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  --local readdatavalid cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1, which is an e_mux
  cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 <= ((cpu_ddr_clock_bridge_s1_readdatavalid_from_sa AND cpu_0_data_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1)) AND NOT cpu_0_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  --cpu_ddr_clock_bridge_s1_writedata mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_writedata <= cpu_0_data_master_writedata;
  --assign cpu_ddr_clock_bridge_s1_endofpacket_from_sa = cpu_ddr_clock_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_ddr_clock_bridge_s1_endofpacket_from_sa <= cpu_ddr_clock_bridge_s1_endofpacket;
  internal_cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 <= ((to_std_logic(((Std_Logic_Vector'(cpu_0_instruction_master_address_to_slave(27 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("0100000000000000000000000000")))) AND (cpu_0_instruction_master_read))) AND cpu_0_instruction_master_read;
  --cpu_0/data_master granted cpu_ddr_clock_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_data_master_granted_slave_cpu_ddr_clock_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_data_master_granted_slave_cpu_ddr_clock_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_data_master_saved_grant_cpu_ddr_clock_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal OR NOT internal_cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_data_master_granted_slave_cpu_ddr_clock_bridge_s1))))));
    end if;

  end process;

  --cpu_0_data_master_continuerequest continued request, which is an e_mux
  cpu_0_data_master_continuerequest <= last_cycle_cpu_0_data_master_granted_slave_cpu_ddr_clock_bridge_s1 AND internal_cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1;
  internal_cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 <= internal_cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 AND NOT ((((cpu_0_instruction_master_read AND (internal_cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register))) OR cpu_0_data_master_arbiterlock));
  --rdv_fifo_for_cpu_0_instruction_master_to_cpu_ddr_clock_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_0_instruction_master_to_cpu_ddr_clock_bridge_s1 : rdv_fifo_for_cpu_0_instruction_master_to_cpu_ddr_clock_bridge_s1_module
    port map(
      data_out => cpu_0_instruction_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1,
      empty => open,
      fifo_contains_ones_n => cpu_0_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1,
      full => open,
      clear_fifo => module_input9,
      clk => clk,
      data_in => internal_cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1,
      read => cpu_ddr_clock_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input10,
      write => module_input11
    );

  module_input9 <= std_logic'('0');
  module_input10 <= std_logic'('0');
  module_input11 <= in_a_read_cycle AND NOT cpu_ddr_clock_bridge_s1_waits_for_read;

  internal_cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register <= NOT cpu_0_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  --local readdatavalid cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1, which is an e_mux
  cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 <= ((cpu_ddr_clock_bridge_s1_readdatavalid_from_sa AND cpu_0_instruction_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1)) AND NOT cpu_0_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  --allow new arb cycle for cpu_ddr_clock_bridge/s1, which is an e_assign
  cpu_ddr_clock_bridge_s1_allow_new_arb_cycle <= NOT cpu_0_data_master_arbiterlock AND NOT cpu_0_instruction_master_arbiterlock;
  --cpu_0/instruction_master assignment into master qualified-requests vector for cpu_ddr_clock_bridge/s1, which is an e_assign
  cpu_ddr_clock_bridge_s1_master_qreq_vector(0) <= internal_cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1;
  --cpu_0/instruction_master grant cpu_ddr_clock_bridge/s1, which is an e_assign
  internal_cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 <= cpu_ddr_clock_bridge_s1_grant_vector(0);
  --cpu_0/instruction_master saved-grant cpu_ddr_clock_bridge/s1, which is an e_assign
  cpu_0_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1 <= cpu_ddr_clock_bridge_s1_arb_winner(0) AND internal_cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  --cpu_0/data_master assignment into master qualified-requests vector for cpu_ddr_clock_bridge/s1, which is an e_assign
  cpu_ddr_clock_bridge_s1_master_qreq_vector(1) <= internal_cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1;
  --cpu_0/data_master grant cpu_ddr_clock_bridge/s1, which is an e_assign
  internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 <= cpu_ddr_clock_bridge_s1_grant_vector(1);
  --cpu_0/data_master saved-grant cpu_ddr_clock_bridge/s1, which is an e_assign
  cpu_0_data_master_saved_grant_cpu_ddr_clock_bridge_s1 <= cpu_ddr_clock_bridge_s1_arb_winner(1) AND internal_cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1;
  --cpu_ddr_clock_bridge/s1 chosen-master double-vector, which is an e_assign
  cpu_ddr_clock_bridge_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((cpu_ddr_clock_bridge_s1_master_qreq_vector & cpu_ddr_clock_bridge_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT cpu_ddr_clock_bridge_s1_master_qreq_vector & NOT cpu_ddr_clock_bridge_s1_master_qreq_vector))) + (std_logic_vector'("000") & (cpu_ddr_clock_bridge_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  cpu_ddr_clock_bridge_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((cpu_ddr_clock_bridge_s1_allow_new_arb_cycle AND or_reduce(cpu_ddr_clock_bridge_s1_grant_vector)))) = '1'), cpu_ddr_clock_bridge_s1_grant_vector, cpu_ddr_clock_bridge_s1_saved_chosen_master_vector);
  --saved cpu_ddr_clock_bridge_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_ddr_clock_bridge_s1_allow_new_arb_cycle) = '1' then 
        cpu_ddr_clock_bridge_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(cpu_ddr_clock_bridge_s1_grant_vector)) = '1'), cpu_ddr_clock_bridge_s1_grant_vector, cpu_ddr_clock_bridge_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  cpu_ddr_clock_bridge_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((cpu_ddr_clock_bridge_s1_chosen_master_double_vector(1) OR cpu_ddr_clock_bridge_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((cpu_ddr_clock_bridge_s1_chosen_master_double_vector(0) OR cpu_ddr_clock_bridge_s1_chosen_master_double_vector(2)))));
  --cpu_ddr_clock_bridge/s1 chosen master rotated left, which is an e_assign
  cpu_ddr_clock_bridge_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(cpu_ddr_clock_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(cpu_ddr_clock_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --cpu_ddr_clock_bridge/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(cpu_ddr_clock_bridge_s1_grant_vector)) = '1' then 
        cpu_ddr_clock_bridge_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(cpu_ddr_clock_bridge_s1_end_xfer) = '1'), cpu_ddr_clock_bridge_s1_chosen_master_rot_left, cpu_ddr_clock_bridge_s1_grant_vector);
      end if;
    end if;

  end process;

  --cpu_ddr_clock_bridge_s1_reset_n assignment, which is an e_assign
  cpu_ddr_clock_bridge_s1_reset_n <= reset_n;
  --cpu_ddr_clock_bridge_s1_firsttransfer first transaction, which is an e_assign
  cpu_ddr_clock_bridge_s1_firsttransfer <= A_WE_StdLogic((std_logic'(cpu_ddr_clock_bridge_s1_begins_xfer) = '1'), cpu_ddr_clock_bridge_s1_unreg_firsttransfer, cpu_ddr_clock_bridge_s1_reg_firsttransfer);
  --cpu_ddr_clock_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  cpu_ddr_clock_bridge_s1_unreg_firsttransfer <= NOT ((cpu_ddr_clock_bridge_s1_slavearbiterlockenable AND cpu_ddr_clock_bridge_s1_any_continuerequest));
  --cpu_ddr_clock_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_ddr_clock_bridge_s1_begins_xfer) = '1' then 
        cpu_ddr_clock_bridge_s1_reg_firsttransfer <= cpu_ddr_clock_bridge_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cpu_ddr_clock_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cpu_ddr_clock_bridge_s1_beginbursttransfer_internal <= cpu_ddr_clock_bridge_s1_begins_xfer;
  --cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal <= cpu_ddr_clock_bridge_s1_begins_xfer AND cpu_ddr_clock_bridge_s1_firsttransfer;
  --cpu_ddr_clock_bridge_s1_read assignment, which is an e_mux
  cpu_ddr_clock_bridge_s1_read <= ((internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 AND cpu_0_data_master_read)) OR ((internal_cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 AND cpu_0_instruction_master_read));
  --cpu_ddr_clock_bridge_s1_write assignment, which is an e_mux
  cpu_ddr_clock_bridge_s1_write <= internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 AND cpu_0_data_master_write;
  shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --cpu_ddr_clock_bridge_s1_address mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1)) = '1'), (A_SRL(shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_0_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 23);
  shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_0_instruction_master <= cpu_0_instruction_master_address_to_slave;
  --slaveid cpu_ddr_clock_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_nativeaddress <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1)) = '1'), (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(cpu_0_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")))), 23);
  --d1_cpu_ddr_clock_bridge_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cpu_ddr_clock_bridge_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cpu_ddr_clock_bridge_s1_end_xfer <= cpu_ddr_clock_bridge_s1_end_xfer;
    end if;

  end process;

  --cpu_ddr_clock_bridge_s1_waits_for_read in a cycle, which is an e_mux
  cpu_ddr_clock_bridge_s1_waits_for_read <= cpu_ddr_clock_bridge_s1_in_a_read_cycle AND internal_cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  --cpu_ddr_clock_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  cpu_ddr_clock_bridge_s1_in_a_read_cycle <= ((internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 AND cpu_0_data_master_read)) OR ((internal_cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 AND cpu_0_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cpu_ddr_clock_bridge_s1_in_a_read_cycle;
  --cpu_ddr_clock_bridge_s1_waits_for_write in a cycle, which is an e_mux
  cpu_ddr_clock_bridge_s1_waits_for_write <= cpu_ddr_clock_bridge_s1_in_a_write_cycle AND internal_cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  --cpu_ddr_clock_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  cpu_ddr_clock_bridge_s1_in_a_write_cycle <= internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cpu_ddr_clock_bridge_s1_in_a_write_cycle;
  wait_for_cpu_ddr_clock_bridge_s1_counter <= std_logic'('0');
  --cpu_ddr_clock_bridge_s1_byteenable byte enable port mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 <= internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 <= internal_cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register <= internal_cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 <= internal_cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 <= internal_cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 <= internal_cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register <= internal_cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 <= internal_cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_s1_waitrequest_from_sa <= internal_cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
--synthesis translate_off
    --cpu_ddr_clock_bridge/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line11 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line11, now);
          write(write_line11, string'(": "));
          write(write_line11, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line11.all);
          deallocate (write_line11);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line12 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_saved_grant_cpu_ddr_clock_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line12, now);
          write(write_line12, string'(": "));
          write(write_line12, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line12.all);
          deallocate (write_line12);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_ddr_clock_bridge_m1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1 : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1_shift_register : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_ddr_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal ddr_sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ddr_sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_ddr_clock_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_latency_counter : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_readdatavalid : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_reset_n : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_waitrequest : OUT STD_LOGIC
              );
end entity cpu_ddr_clock_bridge_m1_arbitrator;


architecture europa of cpu_ddr_clock_bridge_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_read_last_time :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_run :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_write_last_time :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_cpu_ddr_clock_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_cpu_ddr_clock_bridge_m1_waitrequest :  STD_LOGIC;
                signal pre_flush_cpu_ddr_clock_bridge_m1_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 OR NOT cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 OR NOT ((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ddr_sdram_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 OR NOT ((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ddr_sdram_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_ddr_clock_bridge_m1_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_ddr_clock_bridge_m1_address_to_slave <= cpu_ddr_clock_bridge_m1_address(24 DOWNTO 0);
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_cpu_ddr_clock_bridge_m1_readdatavalid <= cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  cpu_ddr_clock_bridge_m1_readdatavalid <= Vector_To_Std_Logic((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_cpu_ddr_clock_bridge_m1_readdatavalid)))));
  --cpu_ddr_clock_bridge/m1 readdata mux, which is an e_mux
  cpu_ddr_clock_bridge_m1_readdata <= ddr_sdram_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_cpu_ddr_clock_bridge_m1_waitrequest <= NOT cpu_ddr_clock_bridge_m1_run;
  --latent max counter, which is an e_assign
  cpu_ddr_clock_bridge_m1_latency_counter <= std_logic'('0');
  --cpu_ddr_clock_bridge_m1_reset_n assignment, which is an e_assign
  cpu_ddr_clock_bridge_m1_reset_n <= reset_n;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_address_to_slave <= internal_cpu_ddr_clock_bridge_m1_address_to_slave;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_waitrequest <= internal_cpu_ddr_clock_bridge_m1_waitrequest;
--synthesis translate_off
    --cpu_ddr_clock_bridge_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_ddr_clock_bridge_m1_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_ddr_clock_bridge_m1_address_last_time <= cpu_ddr_clock_bridge_m1_address;
      end if;

    end process;

    --cpu_ddr_clock_bridge/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpu_ddr_clock_bridge_m1_waitrequest AND ((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write));
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line13 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_ddr_clock_bridge_m1_address /= cpu_ddr_clock_bridge_m1_address_last_time))))) = '1' then 
          write(write_line13, now);
          write(write_line13, string'(": "));
          write(write_line13, string'("cpu_ddr_clock_bridge_m1_address did not heed wait!!!"));
          write(output, write_line13.all);
          deallocate (write_line13);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_ddr_clock_bridge_m1_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        cpu_ddr_clock_bridge_m1_byteenable_last_time <= cpu_ddr_clock_bridge_m1_byteenable;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line14 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_ddr_clock_bridge_m1_byteenable /= cpu_ddr_clock_bridge_m1_byteenable_last_time))))) = '1' then 
          write(write_line14, now);
          write(write_line14, string'(": "));
          write(write_line14, string'("cpu_ddr_clock_bridge_m1_byteenable did not heed wait!!!"));
          write(output, write_line14.all);
          deallocate (write_line14);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_ddr_clock_bridge_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_ddr_clock_bridge_m1_read_last_time <= cpu_ddr_clock_bridge_m1_read;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line15 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_ddr_clock_bridge_m1_read) /= std_logic'(cpu_ddr_clock_bridge_m1_read_last_time)))))) = '1' then 
          write(write_line15, now);
          write(write_line15, string'(": "));
          write(write_line15, string'("cpu_ddr_clock_bridge_m1_read did not heed wait!!!"));
          write(output, write_line15.all);
          deallocate (write_line15);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_ddr_clock_bridge_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_ddr_clock_bridge_m1_write_last_time <= cpu_ddr_clock_bridge_m1_write;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line16 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_ddr_clock_bridge_m1_write) /= std_logic'(cpu_ddr_clock_bridge_m1_write_last_time)))))) = '1' then 
          write(write_line16, now);
          write(write_line16, string'(": "));
          write(write_line16, string'("cpu_ddr_clock_bridge_m1_write did not heed wait!!!"));
          write(output, write_line16.all);
          deallocate (write_line16);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_ddr_clock_bridge_m1_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_ddr_clock_bridge_m1_writedata_last_time <= cpu_ddr_clock_bridge_m1_writedata;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line17 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((cpu_ddr_clock_bridge_m1_writedata /= cpu_ddr_clock_bridge_m1_writedata_last_time)))) AND cpu_ddr_clock_bridge_m1_write)) = '1' then 
          write(write_line17, now);
          write(write_line17, string'(": "));
          write(write_line17, string'("cpu_ddr_clock_bridge_m1_writedata did not heed wait!!!"));
          write(output, write_line17.all);
          deallocate (write_line17);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cpu_ddr_clock_bridge_bridge_arbitrator is 
end entity cpu_ddr_clock_bridge_bridge_arbitrator;


architecture europa of cpu_ddr_clock_bridge_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity dac_ad5308_spi_control_port_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal dac_ad5308_spi_control_port_dataavailable : IN STD_LOGIC;
                 signal dac_ad5308_spi_control_port_endofpacket : IN STD_LOGIC;
                 signal dac_ad5308_spi_control_port_irq : IN STD_LOGIC;
                 signal dac_ad5308_spi_control_port_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal dac_ad5308_spi_control_port_readyfordata : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_3_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal gpib_edm1_clock_3_out_read : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_out_write : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_dac_ad5308_spi_control_port_end_xfer : OUT STD_LOGIC;
                 signal dac_ad5308_spi_control_port_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal dac_ad5308_spi_control_port_chipselect : OUT STD_LOGIC;
                 signal dac_ad5308_spi_control_port_dataavailable_from_sa : OUT STD_LOGIC;
                 signal dac_ad5308_spi_control_port_endofpacket_from_sa : OUT STD_LOGIC;
                 signal dac_ad5308_spi_control_port_irq_from_sa : OUT STD_LOGIC;
                 signal dac_ad5308_spi_control_port_read_n : OUT STD_LOGIC;
                 signal dac_ad5308_spi_control_port_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal dac_ad5308_spi_control_port_readyfordata_from_sa : OUT STD_LOGIC;
                 signal dac_ad5308_spi_control_port_reset_n : OUT STD_LOGIC;
                 signal dac_ad5308_spi_control_port_write_n : OUT STD_LOGIC;
                 signal dac_ad5308_spi_control_port_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_out_read_data_valid_dac_ad5308_spi_control_port : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port : OUT STD_LOGIC
              );
end entity dac_ad5308_spi_control_port_arbitrator;


architecture europa of dac_ad5308_spi_control_port_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_allgrants :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_allow_new_arb_cycle :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_any_bursting_master_saved_grant :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_any_continuerequest :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_arb_counter_enable :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_arb_share_counter :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_arb_share_counter_next_value :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_arb_share_set_values :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_beginbursttransfer_internal :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_begins_xfer :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_end_xfer :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_firsttransfer :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_grant_vector :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_in_a_read_cycle :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_in_a_write_cycle :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_master_qreq_vector :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_non_bursting_master_requests :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_reg_firsttransfer :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_slavearbiterlockenable :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_slavearbiterlockenable2 :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_unreg_firsttransfer :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_waits_for_read :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_waits_for_write :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_dac_ad5308_spi_control_port :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_arbiterlock :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_arbiterlock2 :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_continuerequest :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_saved_grant_dac_ad5308_spi_control_port :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port :  STD_LOGIC;
                signal internal_gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port :  STD_LOGIC;
                signal internal_gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port :  STD_LOGIC;
                signal wait_for_dac_ad5308_spi_control_port_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT dac_ad5308_spi_control_port_end_xfer;
    end if;

  end process;

  dac_ad5308_spi_control_port_begins_xfer <= NOT d1_reasons_to_wait AND (internal_gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port);
  --assign dac_ad5308_spi_control_port_readdata_from_sa = dac_ad5308_spi_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  dac_ad5308_spi_control_port_readdata_from_sa <= dac_ad5308_spi_control_port_readdata;
  internal_gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((gpib_edm1_clock_3_out_read OR gpib_edm1_clock_3_out_write)))))));
  --assign dac_ad5308_spi_control_port_dataavailable_from_sa = dac_ad5308_spi_control_port_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  dac_ad5308_spi_control_port_dataavailable_from_sa <= dac_ad5308_spi_control_port_dataavailable;
  --assign dac_ad5308_spi_control_port_readyfordata_from_sa = dac_ad5308_spi_control_port_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  dac_ad5308_spi_control_port_readyfordata_from_sa <= dac_ad5308_spi_control_port_readyfordata;
  --dac_ad5308_spi_control_port_arb_share_counter set values, which is an e_mux
  dac_ad5308_spi_control_port_arb_share_set_values <= std_logic'('1');
  --dac_ad5308_spi_control_port_non_bursting_master_requests mux, which is an e_mux
  dac_ad5308_spi_control_port_non_bursting_master_requests <= internal_gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port;
  --dac_ad5308_spi_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  dac_ad5308_spi_control_port_any_bursting_master_saved_grant <= std_logic'('0');
  --dac_ad5308_spi_control_port_arb_share_counter_next_value assignment, which is an e_assign
  dac_ad5308_spi_control_port_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(dac_ad5308_spi_control_port_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dac_ad5308_spi_control_port_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(dac_ad5308_spi_control_port_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(dac_ad5308_spi_control_port_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --dac_ad5308_spi_control_port_allgrants all slave grants, which is an e_mux
  dac_ad5308_spi_control_port_allgrants <= dac_ad5308_spi_control_port_grant_vector;
  --dac_ad5308_spi_control_port_end_xfer assignment, which is an e_assign
  dac_ad5308_spi_control_port_end_xfer <= NOT ((dac_ad5308_spi_control_port_waits_for_read OR dac_ad5308_spi_control_port_waits_for_write));
  --end_xfer_arb_share_counter_term_dac_ad5308_spi_control_port arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_dac_ad5308_spi_control_port <= dac_ad5308_spi_control_port_end_xfer AND (((NOT dac_ad5308_spi_control_port_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --dac_ad5308_spi_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  dac_ad5308_spi_control_port_arb_counter_enable <= ((end_xfer_arb_share_counter_term_dac_ad5308_spi_control_port AND dac_ad5308_spi_control_port_allgrants)) OR ((end_xfer_arb_share_counter_term_dac_ad5308_spi_control_port AND NOT dac_ad5308_spi_control_port_non_bursting_master_requests));
  --dac_ad5308_spi_control_port_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dac_ad5308_spi_control_port_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(dac_ad5308_spi_control_port_arb_counter_enable) = '1' then 
        dac_ad5308_spi_control_port_arb_share_counter <= dac_ad5308_spi_control_port_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --dac_ad5308_spi_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dac_ad5308_spi_control_port_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((dac_ad5308_spi_control_port_master_qreq_vector AND end_xfer_arb_share_counter_term_dac_ad5308_spi_control_port)) OR ((end_xfer_arb_share_counter_term_dac_ad5308_spi_control_port AND NOT dac_ad5308_spi_control_port_non_bursting_master_requests)))) = '1' then 
        dac_ad5308_spi_control_port_slavearbiterlockenable <= dac_ad5308_spi_control_port_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_3/out dac_ad5308/spi_control_port arbiterlock, which is an e_assign
  gpib_edm1_clock_3_out_arbiterlock <= dac_ad5308_spi_control_port_slavearbiterlockenable AND gpib_edm1_clock_3_out_continuerequest;
  --dac_ad5308_spi_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  dac_ad5308_spi_control_port_slavearbiterlockenable2 <= dac_ad5308_spi_control_port_arb_share_counter_next_value;
  --gpib_edm1_clock_3/out dac_ad5308/spi_control_port arbiterlock2, which is an e_assign
  gpib_edm1_clock_3_out_arbiterlock2 <= dac_ad5308_spi_control_port_slavearbiterlockenable2 AND gpib_edm1_clock_3_out_continuerequest;
  --dac_ad5308_spi_control_port_any_continuerequest at least one master continues requesting, which is an e_assign
  dac_ad5308_spi_control_port_any_continuerequest <= std_logic'('1');
  --gpib_edm1_clock_3_out_continuerequest continued request, which is an e_assign
  gpib_edm1_clock_3_out_continuerequest <= std_logic'('1');
  internal_gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port <= internal_gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port;
  --dac_ad5308_spi_control_port_writedata mux, which is an e_mux
  dac_ad5308_spi_control_port_writedata <= gpib_edm1_clock_3_out_writedata;
  --assign dac_ad5308_spi_control_port_endofpacket_from_sa = dac_ad5308_spi_control_port_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  dac_ad5308_spi_control_port_endofpacket_from_sa <= dac_ad5308_spi_control_port_endofpacket;
  --master is always granted when requested
  internal_gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port <= internal_gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port;
  --gpib_edm1_clock_3/out saved-grant dac_ad5308/spi_control_port, which is an e_assign
  gpib_edm1_clock_3_out_saved_grant_dac_ad5308_spi_control_port <= internal_gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port;
  --allow new arb cycle for dac_ad5308/spi_control_port, which is an e_assign
  dac_ad5308_spi_control_port_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  dac_ad5308_spi_control_port_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  dac_ad5308_spi_control_port_master_qreq_vector <= std_logic'('1');
  --dac_ad5308_spi_control_port_reset_n assignment, which is an e_assign
  dac_ad5308_spi_control_port_reset_n <= reset_n;
  dac_ad5308_spi_control_port_chipselect <= internal_gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port;
  --dac_ad5308_spi_control_port_firsttransfer first transaction, which is an e_assign
  dac_ad5308_spi_control_port_firsttransfer <= A_WE_StdLogic((std_logic'(dac_ad5308_spi_control_port_begins_xfer) = '1'), dac_ad5308_spi_control_port_unreg_firsttransfer, dac_ad5308_spi_control_port_reg_firsttransfer);
  --dac_ad5308_spi_control_port_unreg_firsttransfer first transaction, which is an e_assign
  dac_ad5308_spi_control_port_unreg_firsttransfer <= NOT ((dac_ad5308_spi_control_port_slavearbiterlockenable AND dac_ad5308_spi_control_port_any_continuerequest));
  --dac_ad5308_spi_control_port_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dac_ad5308_spi_control_port_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(dac_ad5308_spi_control_port_begins_xfer) = '1' then 
        dac_ad5308_spi_control_port_reg_firsttransfer <= dac_ad5308_spi_control_port_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --dac_ad5308_spi_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  dac_ad5308_spi_control_port_beginbursttransfer_internal <= dac_ad5308_spi_control_port_begins_xfer;
  --~dac_ad5308_spi_control_port_read_n assignment, which is an e_mux
  dac_ad5308_spi_control_port_read_n <= NOT ((internal_gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port AND gpib_edm1_clock_3_out_read));
  --~dac_ad5308_spi_control_port_write_n assignment, which is an e_mux
  dac_ad5308_spi_control_port_write_n <= NOT ((internal_gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port AND gpib_edm1_clock_3_out_write));
  --dac_ad5308_spi_control_port_address mux, which is an e_mux
  dac_ad5308_spi_control_port_address <= gpib_edm1_clock_3_out_nativeaddress;
  --d1_dac_ad5308_spi_control_port_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_dac_ad5308_spi_control_port_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_dac_ad5308_spi_control_port_end_xfer <= dac_ad5308_spi_control_port_end_xfer;
    end if;

  end process;

  --dac_ad5308_spi_control_port_waits_for_read in a cycle, which is an e_mux
  dac_ad5308_spi_control_port_waits_for_read <= dac_ad5308_spi_control_port_in_a_read_cycle AND dac_ad5308_spi_control_port_begins_xfer;
  --dac_ad5308_spi_control_port_in_a_read_cycle assignment, which is an e_assign
  dac_ad5308_spi_control_port_in_a_read_cycle <= internal_gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port AND gpib_edm1_clock_3_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= dac_ad5308_spi_control_port_in_a_read_cycle;
  --dac_ad5308_spi_control_port_waits_for_write in a cycle, which is an e_mux
  dac_ad5308_spi_control_port_waits_for_write <= dac_ad5308_spi_control_port_in_a_write_cycle AND dac_ad5308_spi_control_port_begins_xfer;
  --dac_ad5308_spi_control_port_in_a_write_cycle assignment, which is an e_assign
  dac_ad5308_spi_control_port_in_a_write_cycle <= internal_gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port AND gpib_edm1_clock_3_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= dac_ad5308_spi_control_port_in_a_write_cycle;
  wait_for_dac_ad5308_spi_control_port_counter <= std_logic'('0');
  --assign dac_ad5308_spi_control_port_irq_from_sa = dac_ad5308_spi_control_port_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  dac_ad5308_spi_control_port_irq_from_sa <= dac_ad5308_spi_control_port_irq;
  --vhdl renameroo for output signals
  gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port <= internal_gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port;
  --vhdl renameroo for output signals
  gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port <= internal_gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port;
  --vhdl renameroo for output signals
  gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port <= internal_gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port;
--synthesis translate_off
    --dac_ad5308/spi_control_port enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr_sdram_s1_module;


architecture europa of rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ddr_sdram_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ddr_sdram_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ddr_sdram_s1_readdatavalid : IN STD_LOGIC;
                 signal ddr_sdram_s1_resetrequest_n : IN STD_LOGIC;
                 signal ddr_sdram_s1_waitrequest_n : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1 : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 : OUT STD_LOGIC;
                 signal d1_ddr_sdram_s1_end_xfer : OUT STD_LOGIC;
                 signal ddr_sdram_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal ddr_sdram_s1_beginbursttransfer : OUT STD_LOGIC;
                 signal ddr_sdram_s1_burstcount : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal ddr_sdram_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal ddr_sdram_s1_read : OUT STD_LOGIC;
                 signal ddr_sdram_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ddr_sdram_s1_resetrequest_n_from_sa : OUT STD_LOGIC;
                 signal ddr_sdram_s1_waitrequest_n_from_sa : OUT STD_LOGIC;
                 signal ddr_sdram_s1_write : OUT STD_LOGIC;
                 signal ddr_sdram_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity ddr_sdram_s1_arbitrator;


architecture europa of ddr_sdram_s1_arbitrator is
component rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr_sdram_s1_module;

                signal cpu_ddr_clock_bridge_m1_arbiterlock :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_continuerequest :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_rdv_fifo_empty_ddr_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_rdv_fifo_output_from_ddr_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_saved_grant_ddr_sdram_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal ddr_sdram_s1_allgrants :  STD_LOGIC;
                signal ddr_sdram_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal ddr_sdram_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal ddr_sdram_s1_any_continuerequest :  STD_LOGIC;
                signal ddr_sdram_s1_arb_counter_enable :  STD_LOGIC;
                signal ddr_sdram_s1_arb_share_counter :  STD_LOGIC;
                signal ddr_sdram_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal ddr_sdram_s1_arb_share_set_values :  STD_LOGIC;
                signal ddr_sdram_s1_bbt_burstcounter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ddr_sdram_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal ddr_sdram_s1_begins_xfer :  STD_LOGIC;
                signal ddr_sdram_s1_end_xfer :  STD_LOGIC;
                signal ddr_sdram_s1_firsttransfer :  STD_LOGIC;
                signal ddr_sdram_s1_grant_vector :  STD_LOGIC;
                signal ddr_sdram_s1_in_a_read_cycle :  STD_LOGIC;
                signal ddr_sdram_s1_in_a_write_cycle :  STD_LOGIC;
                signal ddr_sdram_s1_master_qreq_vector :  STD_LOGIC;
                signal ddr_sdram_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal ddr_sdram_s1_next_bbt_burstcount :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ddr_sdram_s1_non_bursting_master_requests :  STD_LOGIC;
                signal ddr_sdram_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal ddr_sdram_s1_reg_firsttransfer :  STD_LOGIC;
                signal ddr_sdram_s1_slavearbiterlockenable :  STD_LOGIC;
                signal ddr_sdram_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal ddr_sdram_s1_unreg_firsttransfer :  STD_LOGIC;
                signal ddr_sdram_s1_waits_for_read :  STD_LOGIC;
                signal ddr_sdram_s1_waits_for_write :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_ddr_sdram_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 :  STD_LOGIC;
                signal internal_ddr_sdram_s1_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_ddr_sdram_s1_read :  STD_LOGIC;
                signal internal_ddr_sdram_s1_waitrequest_n_from_sa :  STD_LOGIC;
                signal internal_ddr_sdram_s1_write :  STD_LOGIC;
                signal module_input12 :  STD_LOGIC;
                signal module_input13 :  STD_LOGIC;
                signal module_input14 :  STD_LOGIC;
                signal shifted_address_to_ddr_sdram_s1_from_cpu_ddr_clock_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_ddr_sdram_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT ddr_sdram_s1_end_xfer;
    end if;

  end process;

  ddr_sdram_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1);
  --assign ddr_sdram_s1_readdata_from_sa = ddr_sdram_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  ddr_sdram_s1_readdata_from_sa <= ddr_sdram_s1_readdata;
  internal_cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write)))))));
  --assign ddr_sdram_s1_waitrequest_n_from_sa = ddr_sdram_s1_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_ddr_sdram_s1_waitrequest_n_from_sa <= ddr_sdram_s1_waitrequest_n;
  --assign ddr_sdram_s1_readdatavalid_from_sa = ddr_sdram_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  ddr_sdram_s1_readdatavalid_from_sa <= ddr_sdram_s1_readdatavalid;
  --ddr_sdram_s1_arb_share_counter set values, which is an e_mux
  ddr_sdram_s1_arb_share_set_values <= std_logic'('1');
  --ddr_sdram_s1_non_bursting_master_requests mux, which is an e_mux
  ddr_sdram_s1_non_bursting_master_requests <= internal_cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1;
  --ddr_sdram_s1_any_bursting_master_saved_grant mux, which is an e_mux
  ddr_sdram_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --ddr_sdram_s1_arb_share_counter_next_value assignment, which is an e_assign
  ddr_sdram_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(ddr_sdram_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ddr_sdram_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(ddr_sdram_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ddr_sdram_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --ddr_sdram_s1_allgrants all slave grants, which is an e_mux
  ddr_sdram_s1_allgrants <= ddr_sdram_s1_grant_vector;
  --ddr_sdram_s1_end_xfer assignment, which is an e_assign
  ddr_sdram_s1_end_xfer <= NOT ((ddr_sdram_s1_waits_for_read OR ddr_sdram_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_ddr_sdram_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_ddr_sdram_s1 <= ddr_sdram_s1_end_xfer AND (((NOT ddr_sdram_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --ddr_sdram_s1_arb_share_counter arbitration counter enable, which is an e_assign
  ddr_sdram_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_ddr_sdram_s1 AND ddr_sdram_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_ddr_sdram_s1 AND NOT ddr_sdram_s1_non_bursting_master_requests));
  --ddr_sdram_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ddr_sdram_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(ddr_sdram_s1_arb_counter_enable) = '1' then 
        ddr_sdram_s1_arb_share_counter <= ddr_sdram_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ddr_sdram_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ddr_sdram_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((ddr_sdram_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_ddr_sdram_s1)) OR ((end_xfer_arb_share_counter_term_ddr_sdram_s1 AND NOT ddr_sdram_s1_non_bursting_master_requests)))) = '1' then 
        ddr_sdram_s1_slavearbiterlockenable <= ddr_sdram_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_ddr_clock_bridge/m1 ddr_sdram/s1 arbiterlock, which is an e_assign
  cpu_ddr_clock_bridge_m1_arbiterlock <= ddr_sdram_s1_slavearbiterlockenable AND cpu_ddr_clock_bridge_m1_continuerequest;
  --ddr_sdram_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  ddr_sdram_s1_slavearbiterlockenable2 <= ddr_sdram_s1_arb_share_counter_next_value;
  --cpu_ddr_clock_bridge/m1 ddr_sdram/s1 arbiterlock2, which is an e_assign
  cpu_ddr_clock_bridge_m1_arbiterlock2 <= ddr_sdram_s1_slavearbiterlockenable2 AND cpu_ddr_clock_bridge_m1_continuerequest;
  --ddr_sdram_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  ddr_sdram_s1_any_continuerequest <= std_logic'('1');
  --cpu_ddr_clock_bridge_m1_continuerequest continued request, which is an e_assign
  cpu_ddr_clock_bridge_m1_continuerequest <= std_logic'('1');
  internal_cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 <= internal_cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 AND NOT ((cpu_ddr_clock_bridge_m1_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_m1_latency_counter))))))))));
  --unique name for ddr_sdram_s1_move_on_to_next_transaction, which is an e_assign
  ddr_sdram_s1_move_on_to_next_transaction <= ddr_sdram_s1_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr_sdram_s1 : rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr_sdram_s1_module
    port map(
      data_out => cpu_ddr_clock_bridge_m1_rdv_fifo_output_from_ddr_sdram_s1,
      empty => open,
      fifo_contains_ones_n => cpu_ddr_clock_bridge_m1_rdv_fifo_empty_ddr_sdram_s1,
      full => open,
      clear_fifo => module_input12,
      clk => clk,
      data_in => internal_cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1,
      read => ddr_sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input13,
      write => module_input14
    );

  module_input12 <= std_logic'('0');
  module_input13 <= std_logic'('0');
  module_input14 <= in_a_read_cycle AND NOT ddr_sdram_s1_waits_for_read;

  cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1_shift_register <= NOT cpu_ddr_clock_bridge_m1_rdv_fifo_empty_ddr_sdram_s1;
  --local readdatavalid cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1, which is an e_mux
  cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1 <= ddr_sdram_s1_readdatavalid_from_sa;
  --ddr_sdram_s1_writedata mux, which is an e_mux
  ddr_sdram_s1_writedata <= cpu_ddr_clock_bridge_m1_writedata;
  --master is always granted when requested
  internal_cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 <= internal_cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1;
  --cpu_ddr_clock_bridge/m1 saved-grant ddr_sdram/s1, which is an e_assign
  cpu_ddr_clock_bridge_m1_saved_grant_ddr_sdram_s1 <= internal_cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1;
  --allow new arb cycle for ddr_sdram/s1, which is an e_assign
  ddr_sdram_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  ddr_sdram_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  ddr_sdram_s1_master_qreq_vector <= std_logic'('1');
  --assign ddr_sdram_s1_resetrequest_n_from_sa = ddr_sdram_s1_resetrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  ddr_sdram_s1_resetrequest_n_from_sa <= ddr_sdram_s1_resetrequest_n;
  --ddr_sdram_s1_firsttransfer first transaction, which is an e_assign
  ddr_sdram_s1_firsttransfer <= A_WE_StdLogic((std_logic'(ddr_sdram_s1_begins_xfer) = '1'), ddr_sdram_s1_unreg_firsttransfer, ddr_sdram_s1_reg_firsttransfer);
  --ddr_sdram_s1_unreg_firsttransfer first transaction, which is an e_assign
  ddr_sdram_s1_unreg_firsttransfer <= NOT ((ddr_sdram_s1_slavearbiterlockenable AND ddr_sdram_s1_any_continuerequest));
  --ddr_sdram_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ddr_sdram_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(ddr_sdram_s1_begins_xfer) = '1' then 
        ddr_sdram_s1_reg_firsttransfer <= ddr_sdram_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --ddr_sdram_s1_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  ddr_sdram_s1_next_bbt_burstcount <= A_EXT (A_WE_StdLogicVector((std_logic'((((internal_ddr_sdram_s1_write) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (ddr_sdram_s1_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (internal_ddr_sdram_s1_burstcount)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'((((internal_ddr_sdram_s1_read) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (ddr_sdram_s1_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))))))) = '1'), std_logic_vector'("000000000000000000000000000000000"), (((std_logic_vector'("0000000000000000000000000000000") & (ddr_sdram_s1_bbt_burstcounter)) - std_logic_vector'("000000000000000000000000000000001"))))), 2);
  --ddr_sdram_s1_bbt_burstcounter bbt_burstcounter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ddr_sdram_s1_bbt_burstcounter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(ddr_sdram_s1_begins_xfer) = '1' then 
        ddr_sdram_s1_bbt_burstcounter <= ddr_sdram_s1_next_bbt_burstcount;
      end if;
    end if;

  end process;

  --ddr_sdram_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  ddr_sdram_s1_beginbursttransfer_internal <= ddr_sdram_s1_begins_xfer AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (ddr_sdram_s1_bbt_burstcounter)) = std_logic_vector'("00000000000000000000000000000000"))));
  --ddr_sdram/s1 begin burst transfer to slave, which is an e_assign
  ddr_sdram_s1_beginbursttransfer <= ddr_sdram_s1_beginbursttransfer_internal;
  --ddr_sdram_s1_read assignment, which is an e_mux
  internal_ddr_sdram_s1_read <= internal_cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 AND cpu_ddr_clock_bridge_m1_read;
  --ddr_sdram_s1_write assignment, which is an e_mux
  internal_ddr_sdram_s1_write <= internal_cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 AND cpu_ddr_clock_bridge_m1_write;
  shifted_address_to_ddr_sdram_s1_from_cpu_ddr_clock_bridge_m1 <= cpu_ddr_clock_bridge_m1_address_to_slave;
  --ddr_sdram_s1_address mux, which is an e_mux
  ddr_sdram_s1_address <= A_EXT (A_SRL(shifted_address_to_ddr_sdram_s1_from_cpu_ddr_clock_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 23);
  --d1_ddr_sdram_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_ddr_sdram_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_ddr_sdram_s1_end_xfer <= ddr_sdram_s1_end_xfer;
    end if;

  end process;

  --ddr_sdram_s1_waits_for_read in a cycle, which is an e_mux
  ddr_sdram_s1_waits_for_read <= ddr_sdram_s1_in_a_read_cycle AND NOT internal_ddr_sdram_s1_waitrequest_n_from_sa;
  --ddr_sdram_s1_in_a_read_cycle assignment, which is an e_assign
  ddr_sdram_s1_in_a_read_cycle <= internal_cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 AND cpu_ddr_clock_bridge_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= ddr_sdram_s1_in_a_read_cycle;
  --ddr_sdram_s1_waits_for_write in a cycle, which is an e_mux
  ddr_sdram_s1_waits_for_write <= ddr_sdram_s1_in_a_write_cycle AND NOT internal_ddr_sdram_s1_waitrequest_n_from_sa;
  --ddr_sdram_s1_in_a_write_cycle assignment, which is an e_assign
  ddr_sdram_s1_in_a_write_cycle <= internal_cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 AND cpu_ddr_clock_bridge_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= ddr_sdram_s1_in_a_write_cycle;
  wait_for_ddr_sdram_s1_counter <= std_logic'('0');
  --ddr_sdram_s1_byteenable byte enable port mux, which is an e_mux
  ddr_sdram_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_ddr_clock_bridge_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  internal_ddr_sdram_s1_burstcount <= std_logic_vector'("001");
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 <= internal_cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 <= internal_cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 <= internal_cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1;
  --vhdl renameroo for output signals
  ddr_sdram_s1_burstcount <= internal_ddr_sdram_s1_burstcount;
  --vhdl renameroo for output signals
  ddr_sdram_s1_read <= internal_ddr_sdram_s1_read;
  --vhdl renameroo for output signals
  ddr_sdram_s1_waitrequest_n_from_sa <= internal_ddr_sdram_s1_waitrequest_n_from_sa;
  --vhdl renameroo for output signals
  ddr_sdram_s1_write <= internal_ddr_sdram_s1_write;
--synthesis translate_off
    --ddr_sdram/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_edm1_reset_clk_0_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity gpib_edm1_reset_clk_0_domain_synch_module;


architecture europa of gpib_edm1_reset_clk_0_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_0_data_master_to_flash_ssram_pipeline_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_0_data_master_to_flash_ssram_pipeline_bridge_s1_module;


architecture europa of rdv_fifo_for_cpu_0_data_master_to_flash_ssram_pipeline_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_9;
  empty <= NOT(full_0);
  full_10 <= std_logic'('0');
  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_0_instruction_master_to_flash_ssram_pipeline_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_0_instruction_master_to_flash_ssram_pipeline_bridge_s1_module;


architecture europa of rdv_fifo_for_cpu_0_instruction_master_to_flash_ssram_pipeline_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (4 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_9;
  empty <= NOT(full_0);
  full_10 <= std_logic'('0');
  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 5);
  one_count_minus_one <= A_EXT (((std_logic_vector'("0000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 5);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 5);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity flash_ssram_pipeline_bridge_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_instruction_master_read : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_endofpacket : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_s1_readdatavalid : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal d1_flash_ssram_pipeline_bridge_s1_end_xfer : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_s1_arbiterlock : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_arbiterlock2 : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_burstcount : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_s1_chipselect : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_debugaccess : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_s1_read : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_s1_reset_n : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_write : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity flash_ssram_pipeline_bridge_s1_arbitrator;


architecture europa of flash_ssram_pipeline_bridge_s1_arbitrator is
component rdv_fifo_for_cpu_0_data_master_to_flash_ssram_pipeline_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_0_data_master_to_flash_ssram_pipeline_bridge_s1_module;

component rdv_fifo_for_cpu_0_instruction_master_to_flash_ssram_pipeline_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_0_instruction_master_to_flash_ssram_pipeline_bridge_s1_module;

                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_rdv_fifo_output_from_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_0_instruction_master_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_rdv_fifo_output_from_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_saved_grant_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_allgrants :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_any_continuerequest :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_arb_counter_enable :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_arb_share_counter :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_arb_share_set_values :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_begins_xfer :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_end_xfer :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_firsttransfer :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_in_a_read_cycle :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_in_a_write_cycle :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_non_bursting_master_requests :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_reg_firsttransfer :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_slavearbiterlockenable :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_unreg_firsttransfer :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_waits_for_read :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_flash_ssram_pipeline_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_cpu_0_data_master_granted_slave_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal last_cycle_cpu_0_instruction_master_granted_slave_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal module_input16 :  STD_LOGIC;
                signal module_input17 :  STD_LOGIC;
                signal module_input18 :  STD_LOGIC;
                signal module_input19 :  STD_LOGIC;
                signal module_input20 :  STD_LOGIC;
                signal module_input21 :  STD_LOGIC;
                signal shifted_address_to_flash_ssram_pipeline_bridge_s1_from_cpu_0_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal shifted_address_to_flash_ssram_pipeline_bridge_s1_from_cpu_0_instruction_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_flash_ssram_pipeline_bridge_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT flash_ssram_pipeline_bridge_s1_end_xfer;
    end if;

  end process;

  flash_ssram_pipeline_bridge_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 OR internal_cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1));
  --assign flash_ssram_pipeline_bridge_s1_readdata_from_sa = flash_ssram_pipeline_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  flash_ssram_pipeline_bridge_s1_readdata_from_sa <= flash_ssram_pipeline_bridge_s1_readdata;
  internal_cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(27 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("0110000000000000000000000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign flash_ssram_pipeline_bridge_s1_waitrequest_from_sa = flash_ssram_pipeline_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_flash_ssram_pipeline_bridge_s1_waitrequest_from_sa <= flash_ssram_pipeline_bridge_s1_waitrequest;
  --assign flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa = flash_ssram_pipeline_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa <= flash_ssram_pipeline_bridge_s1_readdatavalid;
  --flash_ssram_pipeline_bridge_s1_arb_share_counter set values, which is an e_mux
  flash_ssram_pipeline_bridge_s1_arb_share_set_values <= std_logic'('1');
  --flash_ssram_pipeline_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  flash_ssram_pipeline_bridge_s1_non_bursting_master_requests <= ((((internal_cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 OR internal_cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1) OR internal_cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1) OR internal_cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1) OR internal_cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1) OR internal_cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1;
  --flash_ssram_pipeline_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  flash_ssram_pipeline_bridge_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(flash_ssram_pipeline_bridge_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(flash_ssram_pipeline_bridge_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(flash_ssram_pipeline_bridge_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(flash_ssram_pipeline_bridge_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --flash_ssram_pipeline_bridge_s1_allgrants all slave grants, which is an e_mux
  flash_ssram_pipeline_bridge_s1_allgrants <= (((((or_reduce(flash_ssram_pipeline_bridge_s1_grant_vector)) OR (or_reduce(flash_ssram_pipeline_bridge_s1_grant_vector))) OR (or_reduce(flash_ssram_pipeline_bridge_s1_grant_vector))) OR (or_reduce(flash_ssram_pipeline_bridge_s1_grant_vector))) OR (or_reduce(flash_ssram_pipeline_bridge_s1_grant_vector))) OR (or_reduce(flash_ssram_pipeline_bridge_s1_grant_vector));
  --flash_ssram_pipeline_bridge_s1_end_xfer assignment, which is an e_assign
  flash_ssram_pipeline_bridge_s1_end_xfer <= NOT ((flash_ssram_pipeline_bridge_s1_waits_for_read OR flash_ssram_pipeline_bridge_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 <= flash_ssram_pipeline_bridge_s1_end_xfer AND (((NOT flash_ssram_pipeline_bridge_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --flash_ssram_pipeline_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  flash_ssram_pipeline_bridge_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 AND flash_ssram_pipeline_bridge_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 AND NOT flash_ssram_pipeline_bridge_s1_non_bursting_master_requests));
  --flash_ssram_pipeline_bridge_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      flash_ssram_pipeline_bridge_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(flash_ssram_pipeline_bridge_s1_arb_counter_enable) = '1' then 
        flash_ssram_pipeline_bridge_s1_arb_share_counter <= flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --flash_ssram_pipeline_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      flash_ssram_pipeline_bridge_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(flash_ssram_pipeline_bridge_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1)) OR ((end_xfer_arb_share_counter_term_flash_ssram_pipeline_bridge_s1 AND NOT flash_ssram_pipeline_bridge_s1_non_bursting_master_requests)))) = '1' then 
        flash_ssram_pipeline_bridge_s1_slavearbiterlockenable <= flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_0/data_master flash_ssram_pipeline_bridge/s1 arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= flash_ssram_pipeline_bridge_s1_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --flash_ssram_pipeline_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  flash_ssram_pipeline_bridge_s1_slavearbiterlockenable2 <= flash_ssram_pipeline_bridge_s1_arb_share_counter_next_value;
  --cpu_0/data_master flash_ssram_pipeline_bridge/s1 arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= flash_ssram_pipeline_bridge_s1_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --cpu_0/instruction_master flash_ssram_pipeline_bridge/s1 arbiterlock, which is an e_assign
  cpu_0_instruction_master_arbiterlock <= flash_ssram_pipeline_bridge_s1_slavearbiterlockenable AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master flash_ssram_pipeline_bridge/s1 arbiterlock2, which is an e_assign
  cpu_0_instruction_master_arbiterlock2 <= flash_ssram_pipeline_bridge_s1_slavearbiterlockenable2 AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master granted flash_ssram_pipeline_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_instruction_master_granted_slave_flash_ssram_pipeline_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_instruction_master_granted_slave_flash_ssram_pipeline_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_instruction_master_saved_grant_flash_ssram_pipeline_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((flash_ssram_pipeline_bridge_s1_arbitration_holdoff_internal OR NOT internal_cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_instruction_master_granted_slave_flash_ssram_pipeline_bridge_s1))))));
    end if;

  end process;

  --cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  cpu_0_instruction_master_continuerequest <= last_cycle_cpu_0_instruction_master_granted_slave_flash_ssram_pipeline_bridge_s1 AND internal_cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1;
  --flash_ssram_pipeline_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  flash_ssram_pipeline_bridge_s1_any_continuerequest <= cpu_0_instruction_master_continuerequest OR cpu_0_data_master_continuerequest;
  internal_cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 <= internal_cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 AND NOT (((((cpu_0_data_master_read AND ((NOT cpu_0_data_master_waitrequest OR (internal_cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register))))) OR (((NOT cpu_0_data_master_waitrequest) AND cpu_0_data_master_write))) OR cpu_0_instruction_master_arbiterlock));
  --unique name for flash_ssram_pipeline_bridge_s1_move_on_to_next_transaction, which is an e_assign
  flash_ssram_pipeline_bridge_s1_move_on_to_next_transaction <= flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_0_data_master_to_flash_ssram_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_0_data_master_to_flash_ssram_pipeline_bridge_s1 : rdv_fifo_for_cpu_0_data_master_to_flash_ssram_pipeline_bridge_s1_module
    port map(
      data_out => cpu_0_data_master_rdv_fifo_output_from_flash_ssram_pipeline_bridge_s1,
      empty => open,
      fifo_contains_ones_n => cpu_0_data_master_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1,
      full => open,
      clear_fifo => module_input16,
      clk => clk,
      data_in => internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1,
      read => flash_ssram_pipeline_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input17,
      write => module_input18
    );

  module_input16 <= std_logic'('0');
  module_input17 <= std_logic'('0');
  module_input18 <= in_a_read_cycle AND NOT flash_ssram_pipeline_bridge_s1_waits_for_read;

  internal_cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register <= NOT cpu_0_data_master_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1;
  --local readdatavalid cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1, which is an e_mux
  cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1 <= ((flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa AND cpu_0_data_master_rdv_fifo_output_from_flash_ssram_pipeline_bridge_s1)) AND NOT cpu_0_data_master_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1;
  --flash_ssram_pipeline_bridge_s1_writedata mux, which is an e_mux
  flash_ssram_pipeline_bridge_s1_writedata <= cpu_0_data_master_writedata;
  --assign flash_ssram_pipeline_bridge_s1_endofpacket_from_sa = flash_ssram_pipeline_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  flash_ssram_pipeline_bridge_s1_endofpacket_from_sa <= flash_ssram_pipeline_bridge_s1_endofpacket;
  internal_cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 <= ((to_std_logic(((Std_Logic_Vector'(cpu_0_instruction_master_address_to_slave(27 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("0110000000000000000000000000")))) AND (cpu_0_instruction_master_read))) AND cpu_0_instruction_master_read;
  --cpu_0/data_master granted flash_ssram_pipeline_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_data_master_granted_slave_flash_ssram_pipeline_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_data_master_granted_slave_flash_ssram_pipeline_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_data_master_saved_grant_flash_ssram_pipeline_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((flash_ssram_pipeline_bridge_s1_arbitration_holdoff_internal OR NOT internal_cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_data_master_granted_slave_flash_ssram_pipeline_bridge_s1))))));
    end if;

  end process;

  --cpu_0_data_master_continuerequest continued request, which is an e_mux
  cpu_0_data_master_continuerequest <= last_cycle_cpu_0_data_master_granted_slave_flash_ssram_pipeline_bridge_s1 AND internal_cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1;
  internal_cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 <= internal_cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 AND NOT ((((cpu_0_instruction_master_read AND (internal_cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register))) OR cpu_0_data_master_arbiterlock));
  --rdv_fifo_for_cpu_0_instruction_master_to_flash_ssram_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_0_instruction_master_to_flash_ssram_pipeline_bridge_s1 : rdv_fifo_for_cpu_0_instruction_master_to_flash_ssram_pipeline_bridge_s1_module
    port map(
      data_out => cpu_0_instruction_master_rdv_fifo_output_from_flash_ssram_pipeline_bridge_s1,
      empty => open,
      fifo_contains_ones_n => cpu_0_instruction_master_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1,
      full => open,
      clear_fifo => module_input19,
      clk => clk,
      data_in => internal_cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1,
      read => flash_ssram_pipeline_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input20,
      write => module_input21
    );

  module_input19 <= std_logic'('0');
  module_input20 <= std_logic'('0');
  module_input21 <= in_a_read_cycle AND NOT flash_ssram_pipeline_bridge_s1_waits_for_read;

  internal_cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register <= NOT cpu_0_instruction_master_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1;
  --local readdatavalid cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1, which is an e_mux
  cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1 <= ((flash_ssram_pipeline_bridge_s1_readdatavalid_from_sa AND cpu_0_instruction_master_rdv_fifo_output_from_flash_ssram_pipeline_bridge_s1)) AND NOT cpu_0_instruction_master_rdv_fifo_empty_flash_ssram_pipeline_bridge_s1;
  --allow new arb cycle for flash_ssram_pipeline_bridge/s1, which is an e_assign
  flash_ssram_pipeline_bridge_s1_allow_new_arb_cycle <= NOT cpu_0_data_master_arbiterlock AND NOT cpu_0_instruction_master_arbiterlock;
  --cpu_0/instruction_master assignment into master qualified-requests vector for flash_ssram_pipeline_bridge/s1, which is an e_assign
  flash_ssram_pipeline_bridge_s1_master_qreq_vector(0) <= internal_cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1;
  --cpu_0/instruction_master grant flash_ssram_pipeline_bridge/s1, which is an e_assign
  internal_cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 <= flash_ssram_pipeline_bridge_s1_grant_vector(0);
  --cpu_0/instruction_master saved-grant flash_ssram_pipeline_bridge/s1, which is an e_assign
  cpu_0_instruction_master_saved_grant_flash_ssram_pipeline_bridge_s1 <= flash_ssram_pipeline_bridge_s1_arb_winner(0) AND internal_cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1;
  --cpu_0/data_master assignment into master qualified-requests vector for flash_ssram_pipeline_bridge/s1, which is an e_assign
  flash_ssram_pipeline_bridge_s1_master_qreq_vector(1) <= internal_cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1;
  --cpu_0/data_master grant flash_ssram_pipeline_bridge/s1, which is an e_assign
  internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 <= flash_ssram_pipeline_bridge_s1_grant_vector(1);
  --cpu_0/data_master saved-grant flash_ssram_pipeline_bridge/s1, which is an e_assign
  cpu_0_data_master_saved_grant_flash_ssram_pipeline_bridge_s1 <= flash_ssram_pipeline_bridge_s1_arb_winner(1) AND internal_cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1;
  --flash_ssram_pipeline_bridge/s1 chosen-master double-vector, which is an e_assign
  flash_ssram_pipeline_bridge_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((flash_ssram_pipeline_bridge_s1_master_qreq_vector & flash_ssram_pipeline_bridge_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT flash_ssram_pipeline_bridge_s1_master_qreq_vector & NOT flash_ssram_pipeline_bridge_s1_master_qreq_vector))) + (std_logic_vector'("000") & (flash_ssram_pipeline_bridge_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  flash_ssram_pipeline_bridge_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((flash_ssram_pipeline_bridge_s1_allow_new_arb_cycle AND or_reduce(flash_ssram_pipeline_bridge_s1_grant_vector)))) = '1'), flash_ssram_pipeline_bridge_s1_grant_vector, flash_ssram_pipeline_bridge_s1_saved_chosen_master_vector);
  --saved flash_ssram_pipeline_bridge_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      flash_ssram_pipeline_bridge_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(flash_ssram_pipeline_bridge_s1_allow_new_arb_cycle) = '1' then 
        flash_ssram_pipeline_bridge_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(flash_ssram_pipeline_bridge_s1_grant_vector)) = '1'), flash_ssram_pipeline_bridge_s1_grant_vector, flash_ssram_pipeline_bridge_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  flash_ssram_pipeline_bridge_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((flash_ssram_pipeline_bridge_s1_chosen_master_double_vector(1) OR flash_ssram_pipeline_bridge_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((flash_ssram_pipeline_bridge_s1_chosen_master_double_vector(0) OR flash_ssram_pipeline_bridge_s1_chosen_master_double_vector(2)))));
  --flash_ssram_pipeline_bridge/s1 chosen master rotated left, which is an e_assign
  flash_ssram_pipeline_bridge_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(flash_ssram_pipeline_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(flash_ssram_pipeline_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --flash_ssram_pipeline_bridge/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      flash_ssram_pipeline_bridge_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(flash_ssram_pipeline_bridge_s1_grant_vector)) = '1' then 
        flash_ssram_pipeline_bridge_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(flash_ssram_pipeline_bridge_s1_end_xfer) = '1'), flash_ssram_pipeline_bridge_s1_chosen_master_rot_left, flash_ssram_pipeline_bridge_s1_grant_vector);
      end if;
    end if;

  end process;

  --flash_ssram_pipeline_bridge_s1_reset_n assignment, which is an e_assign
  flash_ssram_pipeline_bridge_s1_reset_n <= reset_n;
  flash_ssram_pipeline_bridge_s1_chipselect <= internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 OR internal_cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1;
  --flash_ssram_pipeline_bridge_s1_firsttransfer first transaction, which is an e_assign
  flash_ssram_pipeline_bridge_s1_firsttransfer <= A_WE_StdLogic((std_logic'(flash_ssram_pipeline_bridge_s1_begins_xfer) = '1'), flash_ssram_pipeline_bridge_s1_unreg_firsttransfer, flash_ssram_pipeline_bridge_s1_reg_firsttransfer);
  --flash_ssram_pipeline_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  flash_ssram_pipeline_bridge_s1_unreg_firsttransfer <= NOT ((flash_ssram_pipeline_bridge_s1_slavearbiterlockenable AND flash_ssram_pipeline_bridge_s1_any_continuerequest));
  --flash_ssram_pipeline_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      flash_ssram_pipeline_bridge_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(flash_ssram_pipeline_bridge_s1_begins_xfer) = '1' then 
        flash_ssram_pipeline_bridge_s1_reg_firsttransfer <= flash_ssram_pipeline_bridge_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --flash_ssram_pipeline_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  flash_ssram_pipeline_bridge_s1_beginbursttransfer_internal <= flash_ssram_pipeline_bridge_s1_begins_xfer;
  --flash_ssram_pipeline_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  flash_ssram_pipeline_bridge_s1_arbitration_holdoff_internal <= flash_ssram_pipeline_bridge_s1_begins_xfer AND flash_ssram_pipeline_bridge_s1_firsttransfer;
  --flash_ssram_pipeline_bridge_s1_read assignment, which is an e_mux
  flash_ssram_pipeline_bridge_s1_read <= ((internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 AND cpu_0_data_master_read)) OR ((internal_cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 AND cpu_0_instruction_master_read));
  --flash_ssram_pipeline_bridge_s1_write assignment, which is an e_mux
  flash_ssram_pipeline_bridge_s1_write <= internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 AND cpu_0_data_master_write;
  shifted_address_to_flash_ssram_pipeline_bridge_s1_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --flash_ssram_pipeline_bridge_s1_address mux, which is an e_mux
  flash_ssram_pipeline_bridge_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1)) = '1'), (A_SRL(shifted_address_to_flash_ssram_pipeline_bridge_s1_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_flash_ssram_pipeline_bridge_s1_from_cpu_0_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 23);
  shifted_address_to_flash_ssram_pipeline_bridge_s1_from_cpu_0_instruction_master <= cpu_0_instruction_master_address_to_slave;
  --slaveid flash_ssram_pipeline_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  flash_ssram_pipeline_bridge_s1_nativeaddress <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1)) = '1'), (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(cpu_0_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")))), 23);
  --d1_flash_ssram_pipeline_bridge_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_flash_ssram_pipeline_bridge_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_flash_ssram_pipeline_bridge_s1_end_xfer <= flash_ssram_pipeline_bridge_s1_end_xfer;
    end if;

  end process;

  --flash_ssram_pipeline_bridge_s1_waits_for_read in a cycle, which is an e_mux
  flash_ssram_pipeline_bridge_s1_waits_for_read <= flash_ssram_pipeline_bridge_s1_in_a_read_cycle AND internal_flash_ssram_pipeline_bridge_s1_waitrequest_from_sa;
  --flash_ssram_pipeline_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  flash_ssram_pipeline_bridge_s1_in_a_read_cycle <= ((internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 AND cpu_0_data_master_read)) OR ((internal_cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 AND cpu_0_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= flash_ssram_pipeline_bridge_s1_in_a_read_cycle;
  --flash_ssram_pipeline_bridge_s1_waits_for_write in a cycle, which is an e_mux
  flash_ssram_pipeline_bridge_s1_waits_for_write <= flash_ssram_pipeline_bridge_s1_in_a_write_cycle AND internal_flash_ssram_pipeline_bridge_s1_waitrequest_from_sa;
  --flash_ssram_pipeline_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  flash_ssram_pipeline_bridge_s1_in_a_write_cycle <= internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= flash_ssram_pipeline_bridge_s1_in_a_write_cycle;
  wait_for_flash_ssram_pipeline_bridge_s1_counter <= std_logic'('0');
  --flash_ssram_pipeline_bridge_s1_byteenable byte enable port mux, which is an e_mux
  flash_ssram_pipeline_bridge_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  flash_ssram_pipeline_bridge_s1_burstcount <= std_logic'('1');
  --flash_ssram_pipeline_bridge/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  flash_ssram_pipeline_bridge_s1_arbiterlock <= A_WE_StdLogic((std_logic'((cpu_0_data_master_arbiterlock)) = '1'), cpu_0_data_master_arbiterlock, cpu_0_instruction_master_arbiterlock);
  --flash_ssram_pipeline_bridge/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  flash_ssram_pipeline_bridge_s1_arbiterlock2 <= A_WE_StdLogic((std_logic'((cpu_0_data_master_arbiterlock2)) = '1'), cpu_0_data_master_arbiterlock2, cpu_0_instruction_master_arbiterlock2);
  --debugaccess mux, which is an e_mux
  flash_ssram_pipeline_bridge_s1_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 <= internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 <= internal_cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register <= internal_cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 <= internal_cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 <= internal_cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 <= internal_cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register <= internal_cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 <= internal_cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  flash_ssram_pipeline_bridge_s1_waitrequest_from_sa <= internal_flash_ssram_pipeline_bridge_s1_waitrequest_from_sa;
--synthesis translate_off
    --flash_ssram_pipeline_bridge/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line18 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line18, now);
          write(write_line18, string'(": "));
          write(write_line18, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line18.all);
          deallocate (write_line18);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line19 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_saved_grant_flash_ssram_pipeline_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_saved_grant_flash_ssram_pipeline_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line19, now);
          write(write_line19, string'(": "));
          write(write_line19, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line19.all);
          deallocate (write_line19);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity flash_ssram_pipeline_bridge_m1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_pipeline_bridge_before_tristate_s1_end_xfer : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1 : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1_shift_register : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_s1_endofpacket_from_sa : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal flash_ssram_pipeline_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_m1_endofpacket : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_latency_counter : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_m1_readdatavalid : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_waitrequest : OUT STD_LOGIC
              );
end entity flash_ssram_pipeline_bridge_m1_arbitrator;


architecture europa of flash_ssram_pipeline_bridge_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_m1_burstcount_last_time :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_m1_chipselect_last_time :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_read_last_time :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_run :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_write_last_time :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_flash_ssram_pipeline_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_flash_ssram_pipeline_bridge_m1_waitrequest :  STD_LOGIC;
                signal pre_flush_flash_ssram_pipeline_bridge_m1_readdatavalid :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 OR NOT flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 OR NOT flash_ssram_pipeline_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pipeline_bridge_before_tristate_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(flash_ssram_pipeline_bridge_m1_chipselect)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 OR NOT flash_ssram_pipeline_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pipeline_bridge_before_tristate_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(flash_ssram_pipeline_bridge_m1_chipselect)))))))));
  --cascaded wait assignment, which is an e_assign
  flash_ssram_pipeline_bridge_m1_run <= r_2;
  --optimize select-logic by passing only those address bits which matter.
  internal_flash_ssram_pipeline_bridge_m1_address_to_slave <= flash_ssram_pipeline_bridge_m1_address(24 DOWNTO 0);
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_flash_ssram_pipeline_bridge_m1_readdatavalid <= flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  flash_ssram_pipeline_bridge_m1_readdatavalid <= Vector_To_Std_Logic((std_logic_vector'("00000000000000000000000000000000") OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pre_flush_flash_ssram_pipeline_bridge_m1_readdatavalid)))));
  --flash_ssram_pipeline_bridge/m1 readdata mux, which is an e_mux
  flash_ssram_pipeline_bridge_m1_readdata <= pipeline_bridge_before_tristate_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_flash_ssram_pipeline_bridge_m1_waitrequest <= NOT flash_ssram_pipeline_bridge_m1_run;
  --latent max counter, which is an e_assign
  flash_ssram_pipeline_bridge_m1_latency_counter <= std_logic'('0');
  --mux flash_ssram_pipeline_bridge_m1_endofpacket, which is an e_mux
  flash_ssram_pipeline_bridge_m1_endofpacket <= pipeline_bridge_before_tristate_s1_endofpacket_from_sa;
  --vhdl renameroo for output signals
  flash_ssram_pipeline_bridge_m1_address_to_slave <= internal_flash_ssram_pipeline_bridge_m1_address_to_slave;
  --vhdl renameroo for output signals
  flash_ssram_pipeline_bridge_m1_waitrequest <= internal_flash_ssram_pipeline_bridge_m1_waitrequest;
--synthesis translate_off
    --flash_ssram_pipeline_bridge_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        flash_ssram_pipeline_bridge_m1_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        flash_ssram_pipeline_bridge_m1_address_last_time <= flash_ssram_pipeline_bridge_m1_address;
      end if;

    end process;

    --flash_ssram_pipeline_bridge/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_flash_ssram_pipeline_bridge_m1_waitrequest AND flash_ssram_pipeline_bridge_m1_chipselect;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line20 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((flash_ssram_pipeline_bridge_m1_address /= flash_ssram_pipeline_bridge_m1_address_last_time))))) = '1' then 
          write(write_line20, now);
          write(write_line20, string'(": "));
          write(write_line20, string'("flash_ssram_pipeline_bridge_m1_address did not heed wait!!!"));
          write(output, write_line20.all);
          deallocate (write_line20);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_chipselect check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        flash_ssram_pipeline_bridge_m1_chipselect_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        flash_ssram_pipeline_bridge_m1_chipselect_last_time <= flash_ssram_pipeline_bridge_m1_chipselect;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_chipselect matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line21 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(flash_ssram_pipeline_bridge_m1_chipselect) /= std_logic'(flash_ssram_pipeline_bridge_m1_chipselect_last_time)))))) = '1' then 
          write(write_line21, now);
          write(write_line21, string'(": "));
          write(write_line21, string'("flash_ssram_pipeline_bridge_m1_chipselect did not heed wait!!!"));
          write(output, write_line21.all);
          deallocate (write_line21);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        flash_ssram_pipeline_bridge_m1_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        flash_ssram_pipeline_bridge_m1_burstcount_last_time <= flash_ssram_pipeline_bridge_m1_burstcount;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line22 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(flash_ssram_pipeline_bridge_m1_burstcount) /= std_logic'(flash_ssram_pipeline_bridge_m1_burstcount_last_time)))))) = '1' then 
          write(write_line22, now);
          write(write_line22, string'(": "));
          write(write_line22, string'("flash_ssram_pipeline_bridge_m1_burstcount did not heed wait!!!"));
          write(output, write_line22.all);
          deallocate (write_line22);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        flash_ssram_pipeline_bridge_m1_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        flash_ssram_pipeline_bridge_m1_byteenable_last_time <= flash_ssram_pipeline_bridge_m1_byteenable;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line23 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((flash_ssram_pipeline_bridge_m1_byteenable /= flash_ssram_pipeline_bridge_m1_byteenable_last_time))))) = '1' then 
          write(write_line23, now);
          write(write_line23, string'(": "));
          write(write_line23, string'("flash_ssram_pipeline_bridge_m1_byteenable did not heed wait!!!"));
          write(output, write_line23.all);
          deallocate (write_line23);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        flash_ssram_pipeline_bridge_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        flash_ssram_pipeline_bridge_m1_read_last_time <= flash_ssram_pipeline_bridge_m1_read;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line24 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(flash_ssram_pipeline_bridge_m1_read) /= std_logic'(flash_ssram_pipeline_bridge_m1_read_last_time)))))) = '1' then 
          write(write_line24, now);
          write(write_line24, string'(": "));
          write(write_line24, string'("flash_ssram_pipeline_bridge_m1_read did not heed wait!!!"));
          write(output, write_line24.all);
          deallocate (write_line24);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        flash_ssram_pipeline_bridge_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        flash_ssram_pipeline_bridge_m1_write_last_time <= flash_ssram_pipeline_bridge_m1_write;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line25 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(flash_ssram_pipeline_bridge_m1_write) /= std_logic'(flash_ssram_pipeline_bridge_m1_write_last_time)))))) = '1' then 
          write(write_line25, now);
          write(write_line25, string'(": "));
          write(write_line25, string'("flash_ssram_pipeline_bridge_m1_write did not heed wait!!!"));
          write(output, write_line25.all);
          deallocate (write_line25);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        flash_ssram_pipeline_bridge_m1_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        flash_ssram_pipeline_bridge_m1_writedata_last_time <= flash_ssram_pipeline_bridge_m1_writedata;
      end if;

    end process;

    --flash_ssram_pipeline_bridge_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line26 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((flash_ssram_pipeline_bridge_m1_writedata /= flash_ssram_pipeline_bridge_m1_writedata_last_time)))) AND ((flash_ssram_pipeline_bridge_m1_write AND flash_ssram_pipeline_bridge_m1_chipselect)))) = '1' then 
          write(write_line26, now);
          write(write_line26, string'(": "));
          write(write_line26, string'("flash_ssram_pipeline_bridge_m1_writedata did not heed wait!!!"));
          write(output, write_line26.all);
          deallocate (write_line26);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity flash_ssram_pipeline_bridge_bridge_arbitrator is 
end entity flash_ssram_pipeline_bridge_bridge_arbitrator;


architecture europa of flash_ssram_pipeline_bridge_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity flash_ssram_tristate_avalon_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal adsc_n_to_the_ssram : OUT STD_LOGIC;
                 signal bw_n_to_the_ssram : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal bwe_n_to_the_ssram : OUT STD_LOGIC;
                 signal cfi_flash_s1_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal chipenable1_n_to_the_ssram : OUT STD_LOGIC;
                 signal d1_flash_ssram_tristate_avalon_slave_end_xfer : OUT STD_LOGIC;
                 signal flash_ssram_tristate_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal flash_ssram_tristate_data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal incoming_flash_ssram_tristate_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal incoming_flash_ssram_tristate_data_with_Xs_converted_to_0 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal outputenable_n_to_the_ssram : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_granted_ssram_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_requests_ssram_s1 : OUT STD_LOGIC;
                 signal read_n_to_the_cfi_flash : OUT STD_LOGIC;
                 signal reset_n_to_the_ssram : OUT STD_LOGIC;
                 signal select_n_to_the_cfi_flash : OUT STD_LOGIC;
                 signal write_n_to_the_cfi_flash : OUT STD_LOGIC
              );
end entity flash_ssram_tristate_avalon_slave_arbitrator;


architecture europa of flash_ssram_tristate_avalon_slave_arbitrator is
                signal cfi_flash_s1_counter_load_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cfi_flash_s1_in_a_read_cycle :  STD_LOGIC;
                signal cfi_flash_s1_in_a_write_cycle :  STD_LOGIC;
                signal cfi_flash_s1_wait_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cfi_flash_s1_waits_for_read :  STD_LOGIC;
                signal cfi_flash_s1_waits_for_write :  STD_LOGIC;
                signal cfi_flash_s1_with_write_latency :  STD_LOGIC;
                signal d1_in_a_write_cycle :  STD_LOGIC;
                signal d1_outgoing_flash_ssram_tristate_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_flash_ssram_tristate_avalon_slave :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_allgrants :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_any_continuerequest :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_arb_counter_enable :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal flash_ssram_tristate_avalon_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal flash_ssram_tristate_avalon_slave_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal flash_ssram_tristate_avalon_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_begins_xfer :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_end_xfer :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_firsttransfer :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_grant_vector :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_master_qreq_vector :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_non_bursting_master_requests :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_read_pending :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_reg_firsttransfer :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_slavearbiterlockenable :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_unreg_firsttransfer :  STD_LOGIC;
                signal flash_ssram_tristate_avalon_slave_write_pending :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_0_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_10_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_11_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_12_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_13_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_14_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_15_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_1_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_2_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_3_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_4_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_5_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_6_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_7_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_8_is_x :  STD_LOGIC;
                signal incoming_flash_ssram_tristate_data_bit_9_is_x :  STD_LOGIC;
                signal internal_cfi_flash_s1_wait_counter_eq_0 :  STD_LOGIC;
                signal internal_incoming_flash_ssram_tristate_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_before_tristate_m1_granted_ssram_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_before_tristate_m1_requests_ssram_s1 :  STD_LOGIC;
                signal outgoing_flash_ssram_tristate_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_adsc_n_to_the_ssram :  STD_LOGIC;
                signal p1_bw_n_to_the_ssram :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_bwe_n_to_the_ssram :  STD_LOGIC;
                signal p1_chipenable1_n_to_the_ssram :  STD_LOGIC;
                signal p1_flash_ssram_tristate_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal p1_outputenable_n_to_the_ssram :  STD_LOGIC;
                signal p1_pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_read_n_to_the_cfi_flash :  STD_LOGIC;
                signal p1_reset_n_to_the_ssram :  STD_LOGIC;
                signal p1_select_n_to_the_cfi_flash :  STD_LOGIC;
                signal p1_write_n_to_the_cfi_flash :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register_in :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register_in :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_saved_grant_cfi_flash_s1 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_saved_grant_ssram_s1 :  STD_LOGIC;
                signal ssram_s1_in_a_read_cycle :  STD_LOGIC;
                signal ssram_s1_in_a_write_cycle :  STD_LOGIC;
                signal ssram_s1_waits_for_read :  STD_LOGIC;
                signal ssram_s1_waits_for_write :  STD_LOGIC;
                signal ssram_s1_with_write_latency :  STD_LOGIC;
                signal time_to_write :  STD_LOGIC;
                signal wait_for_cfi_flash_s1_counter :  STD_LOGIC;
                signal wait_for_ssram_s1_counter :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of adsc_n_to_the_ssram : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of bw_n_to_the_ssram : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of bwe_n_to_the_ssram : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of chipenable1_n_to_the_ssram : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of d1_in_a_write_cycle : signal is "FAST_OUTPUT_ENABLE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of d1_outgoing_flash_ssram_tristate_data : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of flash_ssram_tristate_address : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of internal_incoming_flash_ssram_tristate_data : signal is "FAST_INPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of outputenable_n_to_the_ssram : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of read_n_to_the_cfi_flash : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of reset_n_to_the_ssram : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of select_n_to_the_cfi_flash : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of write_n_to_the_cfi_flash : signal is "FAST_OUTPUT_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT flash_ssram_tristate_avalon_slave_end_xfer;
    end if;

  end process;

  flash_ssram_tristate_avalon_slave_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 OR internal_pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1));
  internal_pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 <= to_std_logic(((Std_Logic_Vector'(A_ToStdLogicVector(pipeline_bridge_before_tristate_m1_address_to_slave(24)) & std_logic_vector'("000000000000000000000000")) = std_logic_vector'("0000000000000000000000000")))) AND pipeline_bridge_before_tristate_m1_chipselect;
  --~select_n_to_the_cfi_flash of type chipselect to ~p1_select_n_to_the_cfi_flash, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      select_n_to_the_cfi_flash <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      select_n_to_the_cfi_flash <= p1_select_n_to_the_cfi_flash;
    end if;

  end process;

  --~chipenable1_n_to_the_ssram of type chipselect to ~p1_chipenable1_n_to_the_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      chipenable1_n_to_the_ssram <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      chipenable1_n_to_the_ssram <= p1_chipenable1_n_to_the_ssram;
    end if;

  end process;

  flash_ssram_tristate_avalon_slave_write_pending <= std_logic'('0');
  --flash_ssram_tristate/avalon_slave read pending calc, which is an e_assign
  flash_ssram_tristate_avalon_slave_read_pending <= or_reduce(pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register(1 DOWNTO 0));
  --flash_ssram_tristate_avalon_slave_arb_share_counter set values, which is an e_mux
  flash_ssram_tristate_avalon_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000001")), 2);
  --flash_ssram_tristate_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  flash_ssram_tristate_avalon_slave_non_bursting_master_requests <= internal_pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 OR internal_pipeline_bridge_before_tristate_m1_requests_ssram_s1;
  --flash_ssram_tristate_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  flash_ssram_tristate_avalon_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --flash_ssram_tristate_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  flash_ssram_tristate_avalon_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(flash_ssram_tristate_avalon_slave_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (flash_ssram_tristate_avalon_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(flash_ssram_tristate_avalon_slave_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (flash_ssram_tristate_avalon_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --flash_ssram_tristate_avalon_slave_allgrants all slave grants, which is an e_mux
  flash_ssram_tristate_avalon_slave_allgrants <= (flash_ssram_tristate_avalon_slave_grant_vector) OR (flash_ssram_tristate_avalon_slave_grant_vector);
  --flash_ssram_tristate_avalon_slave_end_xfer assignment, which is an e_assign
  flash_ssram_tristate_avalon_slave_end_xfer <= NOT ((((cfi_flash_s1_waits_for_read OR cfi_flash_s1_waits_for_write) OR ssram_s1_waits_for_read) OR ssram_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_flash_ssram_tristate_avalon_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_flash_ssram_tristate_avalon_slave <= flash_ssram_tristate_avalon_slave_end_xfer AND (((NOT flash_ssram_tristate_avalon_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --flash_ssram_tristate_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  flash_ssram_tristate_avalon_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_flash_ssram_tristate_avalon_slave AND flash_ssram_tristate_avalon_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_flash_ssram_tristate_avalon_slave AND NOT flash_ssram_tristate_avalon_slave_non_bursting_master_requests));
  --flash_ssram_tristate_avalon_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      flash_ssram_tristate_avalon_slave_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(flash_ssram_tristate_avalon_slave_arb_counter_enable) = '1' then 
        flash_ssram_tristate_avalon_slave_arb_share_counter <= flash_ssram_tristate_avalon_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --flash_ssram_tristate_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      flash_ssram_tristate_avalon_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((flash_ssram_tristate_avalon_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_flash_ssram_tristate_avalon_slave)) OR ((end_xfer_arb_share_counter_term_flash_ssram_tristate_avalon_slave AND NOT flash_ssram_tristate_avalon_slave_non_bursting_master_requests)))) = '1' then 
        flash_ssram_tristate_avalon_slave_slavearbiterlockenable <= or_reduce(flash_ssram_tristate_avalon_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge_before_tristate/m1 flash_ssram_tristate/avalon_slave arbiterlock, which is an e_assign
  pipeline_bridge_before_tristate_m1_arbiterlock <= flash_ssram_tristate_avalon_slave_slavearbiterlockenable AND pipeline_bridge_before_tristate_m1_continuerequest;
  --flash_ssram_tristate_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  flash_ssram_tristate_avalon_slave_slavearbiterlockenable2 <= or_reduce(flash_ssram_tristate_avalon_slave_arb_share_counter_next_value);
  --pipeline_bridge_before_tristate/m1 flash_ssram_tristate/avalon_slave arbiterlock2, which is an e_assign
  pipeline_bridge_before_tristate_m1_arbiterlock2 <= flash_ssram_tristate_avalon_slave_slavearbiterlockenable2 AND pipeline_bridge_before_tristate_m1_continuerequest;
  --flash_ssram_tristate_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  flash_ssram_tristate_avalon_slave_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_before_tristate_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_before_tristate_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 <= internal_pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 AND NOT ((((((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect)) AND (((flash_ssram_tristate_avalon_slave_write_pending OR (flash_ssram_tristate_avalon_slave_read_pending)) OR to_std_logic(((std_logic_vector'("00000000000000000000000000000010")<(std_logic_vector'("00000000000000000000000000000") & (pipeline_bridge_before_tristate_m1_latency_counter))))))))) OR ((((flash_ssram_tristate_avalon_slave_read_pending OR NOT(or_reduce(internal_pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1)))) AND ((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect))))));
  --pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register_in <= (internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 AND ((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect))) AND NOT cfi_flash_s1_waits_for_read;
  --shift register p1 pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register <= A_EXT ((pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register & A_ToStdLogicVector(pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register_in)), 2);
  --pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register <= p1_pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register;
    end if;

  end process;

  --local readdatavalid pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1, which is an e_mux
  pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1 <= pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1_shift_register(1);
  --flash_ssram_tristate_data register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_incoming_flash_ssram_tristate_data <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      internal_incoming_flash_ssram_tristate_data <= flash_ssram_tristate_data;
    end if;

  end process;

  --cfi_flash_s1_with_write_latency assignment, which is an e_assign
  cfi_flash_s1_with_write_latency <= in_a_write_cycle AND (internal_pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1);
  --time to write the data, which is an e_mux
  time_to_write <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((cfi_flash_s1_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((ssram_s1_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), std_logic_vector'("00000000000000000000000000000000"))));
  --d1_outgoing_flash_ssram_tristate_data register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_outgoing_flash_ssram_tristate_data <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      d1_outgoing_flash_ssram_tristate_data <= outgoing_flash_ssram_tristate_data;
    end if;

  end process;

  --write cycle delayed by 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_in_a_write_cycle <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_in_a_write_cycle <= time_to_write;
    end if;

  end process;

  --d1_outgoing_flash_ssram_tristate_data tristate driver, which is an e_assign
  flash_ssram_tristate_data <= A_WE_StdLogicVector((std_logic'((d1_in_a_write_cycle)) = '1'), d1_outgoing_flash_ssram_tristate_data, A_REP(std_logic'('Z'), 32));
  --outgoing_flash_ssram_tristate_data mux, which is an e_mux
  outgoing_flash_ssram_tristate_data <= A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1)) = '1'), (std_logic_vector'("0000000000000000") & (pipeline_bridge_before_tristate_m1_dbs_write_16)), pipeline_bridge_before_tristate_m1_writedata);
  internal_pipeline_bridge_before_tristate_m1_requests_ssram_s1 <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_before_tristate_m1_address_to_slave(24 DOWNTO 20) & std_logic_vector'("00000000000000000000")) = std_logic_vector'("1000000000000000000000000")))) AND pipeline_bridge_before_tristate_m1_chipselect;
  internal_pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 <= internal_pipeline_bridge_before_tristate_m1_requests_ssram_s1 AND NOT ((((((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect)) AND (((flash_ssram_tristate_avalon_slave_write_pending OR ((flash_ssram_tristate_avalon_slave_read_pending AND NOT((or_reduce(pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register(1 DOWNTO 0))))))) OR to_std_logic(((std_logic_vector'("00000000000000000000000000000100")<(std_logic_vector'("00000000000000000000000000000") & (pipeline_bridge_before_tristate_m1_latency_counter))))))))) OR (((flash_ssram_tristate_avalon_slave_read_pending) AND ((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect))))));
  --pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register_in <= (internal_pipeline_bridge_before_tristate_m1_granted_ssram_s1 AND ((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect))) AND NOT ssram_s1_waits_for_read;
  --shift register p1 pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register <= A_EXT ((pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register & A_ToStdLogicVector(pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register_in)), 4);
  --pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register <= p1_pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register;
    end if;

  end process;

  --local readdatavalid pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1, which is an e_mux
  pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1 <= pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register(3);
  --ssram_s1_with_write_latency assignment, which is an e_assign
  ssram_s1_with_write_latency <= in_a_write_cycle AND (internal_pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1);
  --master is always granted when requested
  internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 <= internal_pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1;
  --pipeline_bridge_before_tristate/m1 saved-grant cfi_flash/s1, which is an e_assign
  pipeline_bridge_before_tristate_m1_saved_grant_cfi_flash_s1 <= internal_pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1;
  --allow new arb cycle for flash_ssram_tristate/avalon_slave, which is an e_assign
  flash_ssram_tristate_avalon_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  flash_ssram_tristate_avalon_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  flash_ssram_tristate_avalon_slave_master_qreq_vector <= std_logic'('1');
  --master is always granted when requested
  internal_pipeline_bridge_before_tristate_m1_granted_ssram_s1 <= internal_pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1;
  --pipeline_bridge_before_tristate/m1 saved-grant ssram/s1, which is an e_assign
  pipeline_bridge_before_tristate_m1_saved_grant_ssram_s1 <= internal_pipeline_bridge_before_tristate_m1_requests_ssram_s1;
  p1_select_n_to_the_cfi_flash <= NOT internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1;
  --flash_ssram_tristate_avalon_slave_firsttransfer first transaction, which is an e_assign
  flash_ssram_tristate_avalon_slave_firsttransfer <= A_WE_StdLogic((std_logic'(flash_ssram_tristate_avalon_slave_begins_xfer) = '1'), flash_ssram_tristate_avalon_slave_unreg_firsttransfer, flash_ssram_tristate_avalon_slave_reg_firsttransfer);
  --flash_ssram_tristate_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  flash_ssram_tristate_avalon_slave_unreg_firsttransfer <= NOT ((flash_ssram_tristate_avalon_slave_slavearbiterlockenable AND flash_ssram_tristate_avalon_slave_any_continuerequest));
  --flash_ssram_tristate_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      flash_ssram_tristate_avalon_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(flash_ssram_tristate_avalon_slave_begins_xfer) = '1' then 
        flash_ssram_tristate_avalon_slave_reg_firsttransfer <= flash_ssram_tristate_avalon_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --flash_ssram_tristate_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  flash_ssram_tristate_avalon_slave_beginbursttransfer_internal <= flash_ssram_tristate_avalon_slave_begins_xfer;
  --~read_n_to_the_cfi_flash of type read to ~p1_read_n_to_the_cfi_flash, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      read_n_to_the_cfi_flash <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      read_n_to_the_cfi_flash <= p1_read_n_to_the_cfi_flash;
    end if;

  end process;

  --~p1_read_n_to_the_cfi_flash assignment, which is an e_mux
  p1_read_n_to_the_cfi_flash <= NOT (((((internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 AND ((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect)))) AND NOT flash_ssram_tristate_avalon_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cfi_flash_s1_wait_counter))<std_logic_vector'("00000000000000000000000000001010"))))));
  --~write_n_to_the_cfi_flash of type write to ~p1_write_n_to_the_cfi_flash, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      write_n_to_the_cfi_flash <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      write_n_to_the_cfi_flash <= p1_write_n_to_the_cfi_flash;
    end if;

  end process;

  --~p1_write_n_to_the_cfi_flash assignment, which is an e_mux
  p1_write_n_to_the_cfi_flash <= NOT ((((((internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 AND ((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect)))) AND NOT flash_ssram_tristate_avalon_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cfi_flash_s1_wait_counter))>=std_logic_vector'("00000000000000000000000000000010"))))) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cfi_flash_s1_wait_counter))<std_logic_vector'("00000000000000000000000000001100"))))));
  --flash_ssram_tristate_address of type address to p1_flash_ssram_tristate_address, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      flash_ssram_tristate_address <= std_logic_vector'("000000000000000000000000");
    elsif clk'event and clk = '1' then
      flash_ssram_tristate_address <= p1_flash_ssram_tristate_address;
    end if;

  end process;

  --p1_flash_ssram_tristate_address mux, which is an e_mux
  p1_flash_ssram_tristate_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1)) = '1'), (Std_Logic_Vector'(A_SRL(pipeline_bridge_before_tristate_m1_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(pipeline_bridge_before_tristate_m1_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0')))), (std_logic_vector'("00") & (pipeline_bridge_before_tristate_m1_address_to_slave))), 24);
  --d1_flash_ssram_tristate_avalon_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_flash_ssram_tristate_avalon_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_flash_ssram_tristate_avalon_slave_end_xfer <= flash_ssram_tristate_avalon_slave_end_xfer;
    end if;

  end process;

  --cfi_flash_s1_waits_for_read in a cycle, which is an e_mux
  cfi_flash_s1_waits_for_read <= cfi_flash_s1_in_a_read_cycle AND wait_for_cfi_flash_s1_counter;
  --cfi_flash_s1_in_a_read_cycle assignment, which is an e_assign
  cfi_flash_s1_in_a_read_cycle <= internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 AND ((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cfi_flash_s1_in_a_read_cycle OR ssram_s1_in_a_read_cycle;
  --cfi_flash_s1_waits_for_write in a cycle, which is an e_mux
  cfi_flash_s1_waits_for_write <= cfi_flash_s1_in_a_write_cycle AND wait_for_cfi_flash_s1_counter;
  --cfi_flash_s1_in_a_write_cycle assignment, which is an e_assign
  cfi_flash_s1_in_a_write_cycle <= internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 AND ((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cfi_flash_s1_in_a_write_cycle OR ssram_s1_in_a_write_cycle;
  internal_cfi_flash_s1_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("0000000000000000000000000000") & (cfi_flash_s1_wait_counter)) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cfi_flash_s1_wait_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      cfi_flash_s1_wait_counter <= cfi_flash_s1_counter_load_value;
    end if;

  end process;

  cfi_flash_s1_counter_load_value <= A_EXT (A_WE_StdLogicVector((std_logic'(((cfi_flash_s1_in_a_read_cycle AND flash_ssram_tristate_avalon_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000001011"), A_WE_StdLogicVector((std_logic'(((cfi_flash_s1_in_a_write_cycle AND flash_ssram_tristate_avalon_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000001101"), A_WE_StdLogicVector((std_logic'((NOT internal_cfi_flash_s1_wait_counter_eq_0)) = '1'), ((std_logic_vector'("00000000000000000000000000000") & (cfi_flash_s1_wait_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000")))), 4);
  wait_for_cfi_flash_s1_counter <= flash_ssram_tristate_avalon_slave_begins_xfer OR NOT internal_cfi_flash_s1_wait_counter_eq_0;
  (pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1_segment_1(1), pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1_segment_1(0), pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1_segment_0(1), pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1_segment_0(0)) <= pipeline_bridge_before_tristate_m1_byteenable;
  internal_pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_before_tristate_m1_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1_segment_0, pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1_segment_1);
  --~adsc_n_to_the_ssram of type begintransfer to ~p1_adsc_n_to_the_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      adsc_n_to_the_ssram <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      adsc_n_to_the_ssram <= p1_adsc_n_to_the_ssram;
    end if;

  end process;

  p1_adsc_n_to_the_ssram <= NOT flash_ssram_tristate_avalon_slave_begins_xfer;
  --~outputenable_n_to_the_ssram of type outputenable to ~p1_outputenable_n_to_the_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      outputenable_n_to_the_ssram <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      outputenable_n_to_the_ssram <= p1_outputenable_n_to_the_ssram;
    end if;

  end process;

  --~p1_outputenable_n_to_the_ssram assignment, which is an e_mux
  p1_outputenable_n_to_the_ssram <= NOT (((or_reduce(pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register(1 DOWNTO 0))) OR ssram_s1_in_a_read_cycle));
  --reset_n_to_the_ssram of type reset_n to p1_reset_n_to_the_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      reset_n_to_the_ssram <= std_logic'('0');
    elsif clk'event and clk = '1' then
      reset_n_to_the_ssram <= p1_reset_n_to_the_ssram;
    end if;

  end process;

  --p1_reset_n_to_the_ssram assignment, which is an e_assign
  p1_reset_n_to_the_ssram <= reset_n;
  p1_chipenable1_n_to_the_ssram <= NOT ((internal_pipeline_bridge_before_tristate_m1_granted_ssram_s1 OR (or_reduce(pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1_shift_register(1 DOWNTO 0)))));
  --~bwe_n_to_the_ssram of type write to ~p1_bwe_n_to_the_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      bwe_n_to_the_ssram <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      bwe_n_to_the_ssram <= p1_bwe_n_to_the_ssram;
    end if;

  end process;

  --~bw_n_to_the_ssram of type byteenable to ~p1_bw_n_to_the_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      bw_n_to_the_ssram <= A_EXT (NOT std_logic_vector'("00000000000000000000000000000000"), 4);
    elsif clk'event and clk = '1' then
      bw_n_to_the_ssram <= p1_bw_n_to_the_ssram;
    end if;

  end process;

  --~p1_bwe_n_to_the_ssram assignment, which is an e_mux
  p1_bwe_n_to_the_ssram <= NOT ((internal_pipeline_bridge_before_tristate_m1_granted_ssram_s1 AND ((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect))));
  --ssram_s1_waits_for_read in a cycle, which is an e_mux
  ssram_s1_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ssram_s1_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --ssram_s1_in_a_read_cycle assignment, which is an e_assign
  ssram_s1_in_a_read_cycle <= internal_pipeline_bridge_before_tristate_m1_granted_ssram_s1 AND ((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect));
  --ssram_s1_waits_for_write in a cycle, which is an e_mux
  ssram_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ssram_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --ssram_s1_in_a_write_cycle assignment, which is an e_assign
  ssram_s1_in_a_write_cycle <= internal_pipeline_bridge_before_tristate_m1_granted_ssram_s1 AND ((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect));
  wait_for_ssram_s1_counter <= std_logic'('0');
  --~p1_bw_n_to_the_ssram byte enable port mux, which is an e_mux
  p1_bw_n_to_the_ssram <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_before_tristate_m1_granted_ssram_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pipeline_bridge_before_tristate_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  --vhdl renameroo for output signals
  cfi_flash_s1_wait_counter_eq_0 <= internal_cfi_flash_s1_wait_counter_eq_0;
  --vhdl renameroo for output signals
  incoming_flash_ssram_tristate_data <= internal_incoming_flash_ssram_tristate_data;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1 <= internal_pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 <= internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_granted_ssram_s1 <= internal_pipeline_bridge_before_tristate_m1_granted_ssram_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 <= internal_pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 <= internal_pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 <= internal_pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_requests_ssram_s1 <= internal_pipeline_bridge_before_tristate_m1_requests_ssram_s1;
--synthesis translate_off
    --incoming_flash_ssram_tristate_data_bit_0_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_0_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(0))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[0] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(0) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_0_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(0));
    --incoming_flash_ssram_tristate_data_bit_1_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_1_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(1))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[1] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(1) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_1_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(1));
    --incoming_flash_ssram_tristate_data_bit_2_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_2_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(2))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[2] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(2) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_2_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(2));
    --incoming_flash_ssram_tristate_data_bit_3_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_3_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(3))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[3] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(3) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_3_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(3));
    --incoming_flash_ssram_tristate_data_bit_4_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_4_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(4))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[4] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(4) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_4_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(4));
    --incoming_flash_ssram_tristate_data_bit_5_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_5_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(5))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[5] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(5) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_5_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(5));
    --incoming_flash_ssram_tristate_data_bit_6_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_6_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(6))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[6] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(6) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_6_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(6));
    --incoming_flash_ssram_tristate_data_bit_7_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_7_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(7))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[7] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(7) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_7_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(7));
    --incoming_flash_ssram_tristate_data_bit_8_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_8_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(8))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[8] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(8) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_8_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(8));
    --incoming_flash_ssram_tristate_data_bit_9_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_9_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(9))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[9] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(9) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_9_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(9));
    --incoming_flash_ssram_tristate_data_bit_10_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_10_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(10))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[10] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(10) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_10_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(10));
    --incoming_flash_ssram_tristate_data_bit_11_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_11_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(11))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[11] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(11) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_11_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(11));
    --incoming_flash_ssram_tristate_data_bit_12_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_12_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(12))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[12] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(12) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_12_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(12));
    --incoming_flash_ssram_tristate_data_bit_13_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_13_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(13))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[13] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(13) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_13_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(13));
    --incoming_flash_ssram_tristate_data_bit_14_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_14_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(14))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[14] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(14) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_14_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(14));
    --incoming_flash_ssram_tristate_data_bit_15_is_x x check, which is an e_assign_is_x
    incoming_flash_ssram_tristate_data_bit_15_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_flash_ssram_tristate_data(15))), '1','0');
    --Crush incoming_flash_ssram_tristate_data_with_Xs_converted_to_0[15] Xs to 0, which is an e_assign
    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(15) <= A_WE_StdLogic((std_logic'(incoming_flash_ssram_tristate_data_bit_15_is_x) = '1'), std_logic'('0'), internal_incoming_flash_ssram_tristate_data(15));
    --cfi_flash/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge_before_tristate/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line27 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_before_tristate_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line27, now);
          write(write_line27, string'(": "));
          write(write_line27, string'("pipeline_bridge_before_tristate/m1 drove 0 on its 'burstcount' port while accessing slave cfi_flash/s1"));
          write(output, write_line27.all);
          deallocate (write_line27);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --ssram/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line28 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pipeline_bridge_before_tristate_m1_granted_ssram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line28, now);
          write(write_line28, string'(": "));
          write(write_line28, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line28.all);
          deallocate (write_line28);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line29 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pipeline_bridge_before_tristate_m1_saved_grant_cfi_flash_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pipeline_bridge_before_tristate_m1_saved_grant_ssram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line29, now);
          write(write_line29, string'(": "));
          write(write_line29, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line29.all);
          deallocate (write_line29);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on
--synthesis read_comments_as_HDL on
--    
--    incoming_flash_ssram_tristate_data_with_Xs_converted_to_0 <= internal_incoming_flash_ssram_tristate_data (15 DOWNTO 0);
--synthesis read_comments_as_HDL off

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity flash_ssram_tristate_bridge_arbitrator is 
end entity flash_ssram_tristate_bridge_arbitrator;


architecture europa of flash_ssram_tristate_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_edm1_clock_0_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpib_edm1_clock_0_in_endofpacket : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_0_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_gpib_edm1_clock_0_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_gpib_edm1_clock_0_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_gpib_edm1_clock_0_in : OUT STD_LOGIC;
                 signal d1_gpib_edm1_clock_0_in_end_xfer : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gpib_edm1_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal gpib_edm1_clock_0_in_read : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_0_in_reset_n : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_in_write : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity gpib_edm1_clock_0_in_arbitrator;


architecture europa of gpib_edm1_clock_0_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_gpib_edm1_clock_0_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gpib_edm1_clock_0_in :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_allgrants :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_allow_new_arb_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_any_continuerequest :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_arb_counter_enable :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_arb_share_counter :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_arb_share_counter_next_value :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_arb_share_set_values :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_beginbursttransfer_internal :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_begins_xfer :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_end_xfer :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_grant_vector :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_in_a_read_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_in_a_write_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_master_qreq_vector :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_non_bursting_master_requests :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_reg_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_slavearbiterlockenable :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_unreg_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_waits_for_read :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_gpib_edm1_clock_0_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_gpib_edm1_clock_0_in :  STD_LOGIC;
                signal internal_gpib_edm1_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal shifted_address_to_gpib_edm1_clock_0_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_gpib_edm1_clock_0_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gpib_edm1_clock_0_in_end_xfer;
    end if;

  end process;

  gpib_edm1_clock_0_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in);
  --assign gpib_edm1_clock_0_in_readdata_from_sa = gpib_edm1_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpib_edm1_clock_0_in_readdata_from_sa <= gpib_edm1_clock_0_in_readdata;
  internal_cpu_0_data_master_requests_gpib_edm1_clock_0_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(27 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1010000000001001000100000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign gpib_edm1_clock_0_in_waitrequest_from_sa = gpib_edm1_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_gpib_edm1_clock_0_in_waitrequest_from_sa <= gpib_edm1_clock_0_in_waitrequest;
  --gpib_edm1_clock_0_in_arb_share_counter set values, which is an e_mux
  gpib_edm1_clock_0_in_arb_share_set_values <= std_logic'('1');
  --gpib_edm1_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  gpib_edm1_clock_0_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_gpib_edm1_clock_0_in;
  --gpib_edm1_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  gpib_edm1_clock_0_in_any_bursting_master_saved_grant <= std_logic'('0');
  --gpib_edm1_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  gpib_edm1_clock_0_in_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gpib_edm1_clock_0_in_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_edm1_clock_0_in_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gpib_edm1_clock_0_in_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_edm1_clock_0_in_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gpib_edm1_clock_0_in_allgrants all slave grants, which is an e_mux
  gpib_edm1_clock_0_in_allgrants <= gpib_edm1_clock_0_in_grant_vector;
  --gpib_edm1_clock_0_in_end_xfer assignment, which is an e_assign
  gpib_edm1_clock_0_in_end_xfer <= NOT ((gpib_edm1_clock_0_in_waits_for_read OR gpib_edm1_clock_0_in_waits_for_write));
  --end_xfer_arb_share_counter_term_gpib_edm1_clock_0_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gpib_edm1_clock_0_in <= gpib_edm1_clock_0_in_end_xfer AND (((NOT gpib_edm1_clock_0_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gpib_edm1_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  gpib_edm1_clock_0_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gpib_edm1_clock_0_in AND gpib_edm1_clock_0_in_allgrants)) OR ((end_xfer_arb_share_counter_term_gpib_edm1_clock_0_in AND NOT gpib_edm1_clock_0_in_non_bursting_master_requests));
  --gpib_edm1_clock_0_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_0_in_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gpib_edm1_clock_0_in_arb_counter_enable) = '1' then 
        gpib_edm1_clock_0_in_arb_share_counter <= gpib_edm1_clock_0_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_0_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gpib_edm1_clock_0_in_master_qreq_vector AND end_xfer_arb_share_counter_term_gpib_edm1_clock_0_in)) OR ((end_xfer_arb_share_counter_term_gpib_edm1_clock_0_in AND NOT gpib_edm1_clock_0_in_non_bursting_master_requests)))) = '1' then 
        gpib_edm1_clock_0_in_slavearbiterlockenable <= gpib_edm1_clock_0_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_0/data_master gpib_edm1_clock_0/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= gpib_edm1_clock_0_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --gpib_edm1_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gpib_edm1_clock_0_in_slavearbiterlockenable2 <= gpib_edm1_clock_0_in_arb_share_counter_next_value;
  --cpu_0/data_master gpib_edm1_clock_0/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= gpib_edm1_clock_0_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --gpib_edm1_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  gpib_edm1_clock_0_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in <= internal_cpu_0_data_master_requests_gpib_edm1_clock_0_in AND NOT ((((cpu_0_data_master_read AND (NOT cpu_0_data_master_waitrequest))) OR (((NOT cpu_0_data_master_waitrequest) AND cpu_0_data_master_write))));
  --gpib_edm1_clock_0_in_writedata mux, which is an e_mux
  gpib_edm1_clock_0_in_writedata <= cpu_0_data_master_writedata (15 DOWNTO 0);
  --assign gpib_edm1_clock_0_in_endofpacket_from_sa = gpib_edm1_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpib_edm1_clock_0_in_endofpacket_from_sa <= gpib_edm1_clock_0_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_gpib_edm1_clock_0_in <= internal_cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in;
  --cpu_0/data_master saved-grant gpib_edm1_clock_0/in, which is an e_assign
  cpu_0_data_master_saved_grant_gpib_edm1_clock_0_in <= internal_cpu_0_data_master_requests_gpib_edm1_clock_0_in;
  --allow new arb cycle for gpib_edm1_clock_0/in, which is an e_assign
  gpib_edm1_clock_0_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gpib_edm1_clock_0_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gpib_edm1_clock_0_in_master_qreq_vector <= std_logic'('1');
  --gpib_edm1_clock_0_in_reset_n assignment, which is an e_assign
  gpib_edm1_clock_0_in_reset_n <= reset_n;
  --gpib_edm1_clock_0_in_firsttransfer first transaction, which is an e_assign
  gpib_edm1_clock_0_in_firsttransfer <= A_WE_StdLogic((std_logic'(gpib_edm1_clock_0_in_begins_xfer) = '1'), gpib_edm1_clock_0_in_unreg_firsttransfer, gpib_edm1_clock_0_in_reg_firsttransfer);
  --gpib_edm1_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  gpib_edm1_clock_0_in_unreg_firsttransfer <= NOT ((gpib_edm1_clock_0_in_slavearbiterlockenable AND gpib_edm1_clock_0_in_any_continuerequest));
  --gpib_edm1_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_0_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gpib_edm1_clock_0_in_begins_xfer) = '1' then 
        gpib_edm1_clock_0_in_reg_firsttransfer <= gpib_edm1_clock_0_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gpib_edm1_clock_0_in_beginbursttransfer_internal <= gpib_edm1_clock_0_in_begins_xfer;
  --gpib_edm1_clock_0_in_read assignment, which is an e_mux
  gpib_edm1_clock_0_in_read <= internal_cpu_0_data_master_granted_gpib_edm1_clock_0_in AND cpu_0_data_master_read;
  --gpib_edm1_clock_0_in_write assignment, which is an e_mux
  gpib_edm1_clock_0_in_write <= internal_cpu_0_data_master_granted_gpib_edm1_clock_0_in AND cpu_0_data_master_write;
  shifted_address_to_gpib_edm1_clock_0_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --gpib_edm1_clock_0_in_address mux, which is an e_mux
  gpib_edm1_clock_0_in_address <= A_EXT (A_SRL(shifted_address_to_gpib_edm1_clock_0_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --slaveid gpib_edm1_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  gpib_edm1_clock_0_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_gpib_edm1_clock_0_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gpib_edm1_clock_0_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gpib_edm1_clock_0_in_end_xfer <= gpib_edm1_clock_0_in_end_xfer;
    end if;

  end process;

  --gpib_edm1_clock_0_in_waits_for_read in a cycle, which is an e_mux
  gpib_edm1_clock_0_in_waits_for_read <= gpib_edm1_clock_0_in_in_a_read_cycle AND internal_gpib_edm1_clock_0_in_waitrequest_from_sa;
  --gpib_edm1_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  gpib_edm1_clock_0_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_gpib_edm1_clock_0_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gpib_edm1_clock_0_in_in_a_read_cycle;
  --gpib_edm1_clock_0_in_waits_for_write in a cycle, which is an e_mux
  gpib_edm1_clock_0_in_waits_for_write <= gpib_edm1_clock_0_in_in_a_write_cycle AND internal_gpib_edm1_clock_0_in_waitrequest_from_sa;
  --gpib_edm1_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  gpib_edm1_clock_0_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_gpib_edm1_clock_0_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gpib_edm1_clock_0_in_in_a_write_cycle;
  wait_for_gpib_edm1_clock_0_in_counter <= std_logic'('0');
  --gpib_edm1_clock_0_in_byteenable byte enable port mux, which is an e_mux
  gpib_edm1_clock_0_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_gpib_edm1_clock_0_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_gpib_edm1_clock_0_in <= internal_cpu_0_data_master_granted_gpib_edm1_clock_0_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in <= internal_cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_gpib_edm1_clock_0_in <= internal_cpu_0_data_master_requests_gpib_edm1_clock_0_in;
  --vhdl renameroo for output signals
  gpib_edm1_clock_0_in_waitrequest_from_sa <= internal_gpib_edm1_clock_0_in_waitrequest_from_sa;
--synthesis translate_off
    --gpib_edm1_clock_0/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity gpib_edm1_clock_0_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_pll_s1_end_xfer : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gpib_edm1_clock_0_out_granted_pll_s1 : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_out_qualified_request_pll_s1 : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_out_read : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_out_read_data_valid_pll_s1 : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_out_requests_pll_s1 : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_out_write : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pll_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal gpib_edm1_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_0_out_reset_n : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_out_waitrequest : OUT STD_LOGIC
              );
end entity gpib_edm1_clock_0_out_arbitrator;


architecture europa of gpib_edm1_clock_0_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_0_out_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_edm1_clock_0_out_read_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_run :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_write_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_gpib_edm1_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_gpib_edm1_clock_0_out_waitrequest :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT gpib_edm1_clock_0_out_qualified_request_pll_s1 OR NOT gpib_edm1_clock_0_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_pll_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_edm1_clock_0_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT gpib_edm1_clock_0_out_qualified_request_pll_s1 OR NOT gpib_edm1_clock_0_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_edm1_clock_0_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  gpib_edm1_clock_0_out_run <= r_2;
  --optimize select-logic by passing only those address bits which matter.
  internal_gpib_edm1_clock_0_out_address_to_slave <= gpib_edm1_clock_0_out_address;
  --gpib_edm1_clock_0/out readdata mux, which is an e_mux
  gpib_edm1_clock_0_out_readdata <= pll_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_gpib_edm1_clock_0_out_waitrequest <= NOT gpib_edm1_clock_0_out_run;
  --gpib_edm1_clock_0_out_reset_n assignment, which is an e_assign
  gpib_edm1_clock_0_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  gpib_edm1_clock_0_out_address_to_slave <= internal_gpib_edm1_clock_0_out_address_to_slave;
  --vhdl renameroo for output signals
  gpib_edm1_clock_0_out_waitrequest <= internal_gpib_edm1_clock_0_out_waitrequest;
--synthesis translate_off
    --gpib_edm1_clock_0_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_0_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_0_out_address_last_time <= gpib_edm1_clock_0_out_address;
      end if;

    end process;

    --gpib_edm1_clock_0/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_gpib_edm1_clock_0_out_waitrequest AND ((gpib_edm1_clock_0_out_read OR gpib_edm1_clock_0_out_write));
      end if;

    end process;

    --gpib_edm1_clock_0_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line30 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_0_out_address /= gpib_edm1_clock_0_out_address_last_time))))) = '1' then 
          write(write_line30, now);
          write(write_line30, string'(": "));
          write(write_line30, string'("gpib_edm1_clock_0_out_address did not heed wait!!!"));
          write(output, write_line30.all);
          deallocate (write_line30);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_0_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_0_out_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_0_out_byteenable_last_time <= gpib_edm1_clock_0_out_byteenable;
      end if;

    end process;

    --gpib_edm1_clock_0_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line31 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_0_out_byteenable /= gpib_edm1_clock_0_out_byteenable_last_time))))) = '1' then 
          write(write_line31, now);
          write(write_line31, string'(": "));
          write(write_line31, string'("gpib_edm1_clock_0_out_byteenable did not heed wait!!!"));
          write(output, write_line31.all);
          deallocate (write_line31);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_0_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_0_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_0_out_read_last_time <= gpib_edm1_clock_0_out_read;
      end if;

    end process;

    --gpib_edm1_clock_0_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line32 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(gpib_edm1_clock_0_out_read) /= std_logic'(gpib_edm1_clock_0_out_read_last_time)))))) = '1' then 
          write(write_line32, now);
          write(write_line32, string'(": "));
          write(write_line32, string'("gpib_edm1_clock_0_out_read did not heed wait!!!"));
          write(output, write_line32.all);
          deallocate (write_line32);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_0_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_0_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_0_out_write_last_time <= gpib_edm1_clock_0_out_write;
      end if;

    end process;

    --gpib_edm1_clock_0_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line33 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(gpib_edm1_clock_0_out_write) /= std_logic'(gpib_edm1_clock_0_out_write_last_time)))))) = '1' then 
          write(write_line33, now);
          write(write_line33, string'(": "));
          write(write_line33, string'("gpib_edm1_clock_0_out_write did not heed wait!!!"));
          write(output, write_line33.all);
          deallocate (write_line33);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_0_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_0_out_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_0_out_writedata_last_time <= gpib_edm1_clock_0_out_writedata;
      end if;

    end process;

    --gpib_edm1_clock_0_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line34 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_0_out_writedata /= gpib_edm1_clock_0_out_writedata_last_time)))) AND gpib_edm1_clock_0_out_write)) = '1' then 
          write(write_line34, now);
          write(write_line34, string'(": "));
          write(write_line34, string'("gpib_edm1_clock_0_out_writedata did not heed wait!!!"));
          write(output, write_line34.all);
          deallocate (write_line34);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_edm1_clock_1_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpib_edm1_clock_1_in_endofpacket : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpib_edm1_clock_1_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_gpib_edm1_clock_1_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_gpib_edm1_clock_1_in : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_gpib_edm1_clock_1_in : OUT STD_LOGIC;
                 signal d1_gpib_edm1_clock_1_in_end_xfer : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_in_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gpib_edm1_clock_1_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_1_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_in_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal gpib_edm1_clock_1_in_read : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpib_edm1_clock_1_in_reset_n : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_in_write : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity gpib_edm1_clock_1_in_arbitrator;


architecture europa of gpib_edm1_clock_1_in_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_gpib_edm1_clock_1_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gpib_edm1_clock_1_in :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_allgrants :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_allow_new_arb_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_any_continuerequest :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_arb_counter_enable :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_arb_share_counter :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_arb_share_counter_next_value :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_arb_share_set_values :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_beginbursttransfer_internal :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_begins_xfer :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_end_xfer :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_grant_vector :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_in_a_read_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_in_a_write_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_master_qreq_vector :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_non_bursting_master_requests :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_reg_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_slavearbiterlockenable :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_unreg_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_waits_for_read :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_gpib_edm1_clock_1_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_gpib_edm1_clock_1_in :  STD_LOGIC;
                signal internal_gpib_edm1_clock_1_in_waitrequest_from_sa :  STD_LOGIC;
                signal shifted_address_to_gpib_edm1_clock_1_in_from_cpu_0_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_gpib_edm1_clock_1_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gpib_edm1_clock_1_in_end_xfer;
    end if;

  end process;

  gpib_edm1_clock_1_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in);
  --assign gpib_edm1_clock_1_in_readdata_from_sa = gpib_edm1_clock_1_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpib_edm1_clock_1_in_readdata_from_sa <= gpib_edm1_clock_1_in_readdata;
  internal_cpu_0_data_master_requests_gpib_edm1_clock_1_in <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(27 DOWNTO 8) & std_logic_vector'("00000000")) = std_logic_vector'("1010000000001001000000000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --assign gpib_edm1_clock_1_in_waitrequest_from_sa = gpib_edm1_clock_1_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_gpib_edm1_clock_1_in_waitrequest_from_sa <= gpib_edm1_clock_1_in_waitrequest;
  --gpib_edm1_clock_1_in_arb_share_counter set values, which is an e_mux
  gpib_edm1_clock_1_in_arb_share_set_values <= std_logic'('1');
  --gpib_edm1_clock_1_in_non_bursting_master_requests mux, which is an e_mux
  gpib_edm1_clock_1_in_non_bursting_master_requests <= internal_cpu_0_data_master_requests_gpib_edm1_clock_1_in;
  --gpib_edm1_clock_1_in_any_bursting_master_saved_grant mux, which is an e_mux
  gpib_edm1_clock_1_in_any_bursting_master_saved_grant <= std_logic'('0');
  --gpib_edm1_clock_1_in_arb_share_counter_next_value assignment, which is an e_assign
  gpib_edm1_clock_1_in_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gpib_edm1_clock_1_in_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_edm1_clock_1_in_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gpib_edm1_clock_1_in_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_edm1_clock_1_in_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gpib_edm1_clock_1_in_allgrants all slave grants, which is an e_mux
  gpib_edm1_clock_1_in_allgrants <= gpib_edm1_clock_1_in_grant_vector;
  --gpib_edm1_clock_1_in_end_xfer assignment, which is an e_assign
  gpib_edm1_clock_1_in_end_xfer <= NOT ((gpib_edm1_clock_1_in_waits_for_read OR gpib_edm1_clock_1_in_waits_for_write));
  --end_xfer_arb_share_counter_term_gpib_edm1_clock_1_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gpib_edm1_clock_1_in <= gpib_edm1_clock_1_in_end_xfer AND (((NOT gpib_edm1_clock_1_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gpib_edm1_clock_1_in_arb_share_counter arbitration counter enable, which is an e_assign
  gpib_edm1_clock_1_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gpib_edm1_clock_1_in AND gpib_edm1_clock_1_in_allgrants)) OR ((end_xfer_arb_share_counter_term_gpib_edm1_clock_1_in AND NOT gpib_edm1_clock_1_in_non_bursting_master_requests));
  --gpib_edm1_clock_1_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_1_in_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gpib_edm1_clock_1_in_arb_counter_enable) = '1' then 
        gpib_edm1_clock_1_in_arb_share_counter <= gpib_edm1_clock_1_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_1_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_1_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gpib_edm1_clock_1_in_master_qreq_vector AND end_xfer_arb_share_counter_term_gpib_edm1_clock_1_in)) OR ((end_xfer_arb_share_counter_term_gpib_edm1_clock_1_in AND NOT gpib_edm1_clock_1_in_non_bursting_master_requests)))) = '1' then 
        gpib_edm1_clock_1_in_slavearbiterlockenable <= gpib_edm1_clock_1_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_0/data_master gpib_edm1_clock_1/in arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= gpib_edm1_clock_1_in_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --gpib_edm1_clock_1_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gpib_edm1_clock_1_in_slavearbiterlockenable2 <= gpib_edm1_clock_1_in_arb_share_counter_next_value;
  --cpu_0/data_master gpib_edm1_clock_1/in arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= gpib_edm1_clock_1_in_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --gpib_edm1_clock_1_in_any_continuerequest at least one master continues requesting, which is an e_assign
  gpib_edm1_clock_1_in_any_continuerequest <= std_logic'('1');
  --cpu_0_data_master_continuerequest continued request, which is an e_assign
  cpu_0_data_master_continuerequest <= std_logic'('1');
  internal_cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in <= internal_cpu_0_data_master_requests_gpib_edm1_clock_1_in AND NOT ((((cpu_0_data_master_read AND (NOT cpu_0_data_master_waitrequest))) OR (((NOT cpu_0_data_master_waitrequest) AND cpu_0_data_master_write))));
  --gpib_edm1_clock_1_in_writedata mux, which is an e_mux
  gpib_edm1_clock_1_in_writedata <= cpu_0_data_master_writedata;
  --assign gpib_edm1_clock_1_in_endofpacket_from_sa = gpib_edm1_clock_1_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpib_edm1_clock_1_in_endofpacket_from_sa <= gpib_edm1_clock_1_in_endofpacket;
  --master is always granted when requested
  internal_cpu_0_data_master_granted_gpib_edm1_clock_1_in <= internal_cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in;
  --cpu_0/data_master saved-grant gpib_edm1_clock_1/in, which is an e_assign
  cpu_0_data_master_saved_grant_gpib_edm1_clock_1_in <= internal_cpu_0_data_master_requests_gpib_edm1_clock_1_in;
  --allow new arb cycle for gpib_edm1_clock_1/in, which is an e_assign
  gpib_edm1_clock_1_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gpib_edm1_clock_1_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gpib_edm1_clock_1_in_master_qreq_vector <= std_logic'('1');
  --gpib_edm1_clock_1_in_reset_n assignment, which is an e_assign
  gpib_edm1_clock_1_in_reset_n <= reset_n;
  --gpib_edm1_clock_1_in_firsttransfer first transaction, which is an e_assign
  gpib_edm1_clock_1_in_firsttransfer <= A_WE_StdLogic((std_logic'(gpib_edm1_clock_1_in_begins_xfer) = '1'), gpib_edm1_clock_1_in_unreg_firsttransfer, gpib_edm1_clock_1_in_reg_firsttransfer);
  --gpib_edm1_clock_1_in_unreg_firsttransfer first transaction, which is an e_assign
  gpib_edm1_clock_1_in_unreg_firsttransfer <= NOT ((gpib_edm1_clock_1_in_slavearbiterlockenable AND gpib_edm1_clock_1_in_any_continuerequest));
  --gpib_edm1_clock_1_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_1_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gpib_edm1_clock_1_in_begins_xfer) = '1' then 
        gpib_edm1_clock_1_in_reg_firsttransfer <= gpib_edm1_clock_1_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_1_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gpib_edm1_clock_1_in_beginbursttransfer_internal <= gpib_edm1_clock_1_in_begins_xfer;
  --gpib_edm1_clock_1_in_read assignment, which is an e_mux
  gpib_edm1_clock_1_in_read <= internal_cpu_0_data_master_granted_gpib_edm1_clock_1_in AND cpu_0_data_master_read;
  --gpib_edm1_clock_1_in_write assignment, which is an e_mux
  gpib_edm1_clock_1_in_write <= internal_cpu_0_data_master_granted_gpib_edm1_clock_1_in AND cpu_0_data_master_write;
  shifted_address_to_gpib_edm1_clock_1_in_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --gpib_edm1_clock_1_in_address mux, which is an e_mux
  gpib_edm1_clock_1_in_address <= A_EXT (A_SRL(shifted_address_to_gpib_edm1_clock_1_in_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010")), 8);
  --slaveid gpib_edm1_clock_1_in_nativeaddress nativeaddress mux, which is an e_mux
  gpib_edm1_clock_1_in_nativeaddress <= A_EXT (A_SRL(cpu_0_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 6);
  --d1_gpib_edm1_clock_1_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gpib_edm1_clock_1_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gpib_edm1_clock_1_in_end_xfer <= gpib_edm1_clock_1_in_end_xfer;
    end if;

  end process;

  --gpib_edm1_clock_1_in_waits_for_read in a cycle, which is an e_mux
  gpib_edm1_clock_1_in_waits_for_read <= gpib_edm1_clock_1_in_in_a_read_cycle AND internal_gpib_edm1_clock_1_in_waitrequest_from_sa;
  --gpib_edm1_clock_1_in_in_a_read_cycle assignment, which is an e_assign
  gpib_edm1_clock_1_in_in_a_read_cycle <= internal_cpu_0_data_master_granted_gpib_edm1_clock_1_in AND cpu_0_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gpib_edm1_clock_1_in_in_a_read_cycle;
  --gpib_edm1_clock_1_in_waits_for_write in a cycle, which is an e_mux
  gpib_edm1_clock_1_in_waits_for_write <= gpib_edm1_clock_1_in_in_a_write_cycle AND internal_gpib_edm1_clock_1_in_waitrequest_from_sa;
  --gpib_edm1_clock_1_in_in_a_write_cycle assignment, which is an e_assign
  gpib_edm1_clock_1_in_in_a_write_cycle <= internal_cpu_0_data_master_granted_gpib_edm1_clock_1_in AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gpib_edm1_clock_1_in_in_a_write_cycle;
  wait_for_gpib_edm1_clock_1_in_counter <= std_logic'('0');
  --gpib_edm1_clock_1_in_byteenable byte enable port mux, which is an e_mux
  gpib_edm1_clock_1_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_gpib_edm1_clock_1_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_gpib_edm1_clock_1_in <= internal_cpu_0_data_master_granted_gpib_edm1_clock_1_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in <= internal_cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_gpib_edm1_clock_1_in <= internal_cpu_0_data_master_requests_gpib_edm1_clock_1_in;
  --vhdl renameroo for output signals
  gpib_edm1_clock_1_in_waitrequest_from_sa <= internal_gpib_edm1_clock_1_in_waitrequest_from_sa;
--synthesis translate_off
    --gpib_edm1_clock_1/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity gpib_edm1_clock_1_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_remote_update_cycloneiii_1_s1_end_xfer : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_out_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gpib_edm1_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_out_read : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1 : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_out_write : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal remote_update_cycloneiii_1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal remote_update_cycloneiii_1_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal gpib_edm1_clock_1_out_address_to_slave : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gpib_edm1_clock_1_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpib_edm1_clock_1_out_reset_n : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_out_waitrequest : OUT STD_LOGIC
              );
end entity gpib_edm1_clock_1_out_arbitrator;


architecture europa of gpib_edm1_clock_1_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_address_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpib_edm1_clock_1_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_1_out_read_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_run :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_write_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_gpib_edm1_clock_1_out_address_to_slave :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_gpib_edm1_clock_1_out_waitrequest :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 OR gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1) OR NOT gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 OR NOT gpib_edm1_clock_1_out_read) OR ((gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1 AND gpib_edm1_clock_1_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 OR NOT ((gpib_edm1_clock_1_out_read OR gpib_edm1_clock_1_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT remote_update_cycloneiii_1_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((gpib_edm1_clock_1_out_read OR gpib_edm1_clock_1_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  gpib_edm1_clock_1_out_run <= r_2;
  --optimize select-logic by passing only those address bits which matter.
  internal_gpib_edm1_clock_1_out_address_to_slave <= gpib_edm1_clock_1_out_address;
  --gpib_edm1_clock_1/out readdata mux, which is an e_mux
  gpib_edm1_clock_1_out_readdata <= remote_update_cycloneiii_1_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_gpib_edm1_clock_1_out_waitrequest <= NOT gpib_edm1_clock_1_out_run;
  --gpib_edm1_clock_1_out_reset_n assignment, which is an e_assign
  gpib_edm1_clock_1_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  gpib_edm1_clock_1_out_address_to_slave <= internal_gpib_edm1_clock_1_out_address_to_slave;
  --vhdl renameroo for output signals
  gpib_edm1_clock_1_out_waitrequest <= internal_gpib_edm1_clock_1_out_waitrequest;
--synthesis translate_off
    --gpib_edm1_clock_1_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_1_out_address_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_1_out_address_last_time <= gpib_edm1_clock_1_out_address;
      end if;

    end process;

    --gpib_edm1_clock_1/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_gpib_edm1_clock_1_out_waitrequest AND ((gpib_edm1_clock_1_out_read OR gpib_edm1_clock_1_out_write));
      end if;

    end process;

    --gpib_edm1_clock_1_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line35 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_1_out_address /= gpib_edm1_clock_1_out_address_last_time))))) = '1' then 
          write(write_line35, now);
          write(write_line35, string'(": "));
          write(write_line35, string'("gpib_edm1_clock_1_out_address did not heed wait!!!"));
          write(output, write_line35.all);
          deallocate (write_line35);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_1_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_1_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_1_out_byteenable_last_time <= gpib_edm1_clock_1_out_byteenable;
      end if;

    end process;

    --gpib_edm1_clock_1_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line36 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_1_out_byteenable /= gpib_edm1_clock_1_out_byteenable_last_time))))) = '1' then 
          write(write_line36, now);
          write(write_line36, string'(": "));
          write(write_line36, string'("gpib_edm1_clock_1_out_byteenable did not heed wait!!!"));
          write(output, write_line36.all);
          deallocate (write_line36);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_1_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_1_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_1_out_read_last_time <= gpib_edm1_clock_1_out_read;
      end if;

    end process;

    --gpib_edm1_clock_1_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line37 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(gpib_edm1_clock_1_out_read) /= std_logic'(gpib_edm1_clock_1_out_read_last_time)))))) = '1' then 
          write(write_line37, now);
          write(write_line37, string'(": "));
          write(write_line37, string'("gpib_edm1_clock_1_out_read did not heed wait!!!"));
          write(output, write_line37.all);
          deallocate (write_line37);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_1_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_1_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_1_out_write_last_time <= gpib_edm1_clock_1_out_write;
      end if;

    end process;

    --gpib_edm1_clock_1_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line38 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(gpib_edm1_clock_1_out_write) /= std_logic'(gpib_edm1_clock_1_out_write_last_time)))))) = '1' then 
          write(write_line38, now);
          write(write_line38, string'(": "));
          write(write_line38, string'("gpib_edm1_clock_1_out_write did not heed wait!!!"));
          write(output, write_line38.all);
          deallocate (write_line38);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_1_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_1_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_1_out_writedata_last_time <= gpib_edm1_clock_1_out_writedata;
      end if;

    end process;

    --gpib_edm1_clock_1_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line39 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_1_out_writedata /= gpib_edm1_clock_1_out_writedata_last_time)))) AND gpib_edm1_clock_1_out_write)) = '1' then 
          write(write_line39, now);
          write(write_line39, string'(": "));
          write(write_line39, string'("gpib_edm1_clock_1_out_writedata did not heed wait!!!"));
          write(output, write_line39.all);
          deallocate (write_line39);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_edm1_clock_2_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpib_edm1_clock_2_in_endofpacket : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_2_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_m1_granted_gpib_edm1_clock_2_in : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_gpib_edm1_clock_2_in : OUT STD_LOGIC;
                 signal d1_gpib_edm1_clock_2_in_end_xfer : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_2_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gpib_edm1_clock_2_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal gpib_edm1_clock_2_in_read : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_2_in_reset_n : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_in_write : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity gpib_edm1_clock_2_in_arbitrator;


architecture europa of gpib_edm1_clock_2_in_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_gpib_edm1_clock_2_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gpib_edm1_clock_2_in :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_allgrants :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_allow_new_arb_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_any_continuerequest :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_arb_counter_enable :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_arb_share_counter :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_arb_share_counter_next_value :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_arb_share_set_values :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_beginbursttransfer_internal :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_begins_xfer :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_end_xfer :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_grant_vector :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_in_a_read_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_in_a_write_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_master_qreq_vector :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_non_bursting_master_requests :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_reg_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_slavearbiterlockenable :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_unreg_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_waits_for_read :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_gpib_edm1_clock_2_in :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_gpib_edm1_clock_2_in :  STD_LOGIC;
                signal internal_gpib_edm1_clock_2_in_waitrequest_from_sa :  STD_LOGIC;
                signal wait_for_gpib_edm1_clock_2_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gpib_edm1_clock_2_in_end_xfer;
    end if;

  end process;

  gpib_edm1_clock_2_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in);
  --assign gpib_edm1_clock_2_in_readdata_from_sa = gpib_edm1_clock_2_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpib_edm1_clock_2_in_readdata_from_sa <= gpib_edm1_clock_2_in_readdata;
  internal_clock_crossing_0_m1_requests_gpib_edm1_clock_2_in <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(7 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("01100000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --assign gpib_edm1_clock_2_in_waitrequest_from_sa = gpib_edm1_clock_2_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_gpib_edm1_clock_2_in_waitrequest_from_sa <= gpib_edm1_clock_2_in_waitrequest;
  --gpib_edm1_clock_2_in_arb_share_counter set values, which is an e_mux
  gpib_edm1_clock_2_in_arb_share_set_values <= std_logic'('1');
  --gpib_edm1_clock_2_in_non_bursting_master_requests mux, which is an e_mux
  gpib_edm1_clock_2_in_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_gpib_edm1_clock_2_in;
  --gpib_edm1_clock_2_in_any_bursting_master_saved_grant mux, which is an e_mux
  gpib_edm1_clock_2_in_any_bursting_master_saved_grant <= std_logic'('0');
  --gpib_edm1_clock_2_in_arb_share_counter_next_value assignment, which is an e_assign
  gpib_edm1_clock_2_in_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gpib_edm1_clock_2_in_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_edm1_clock_2_in_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gpib_edm1_clock_2_in_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_edm1_clock_2_in_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gpib_edm1_clock_2_in_allgrants all slave grants, which is an e_mux
  gpib_edm1_clock_2_in_allgrants <= gpib_edm1_clock_2_in_grant_vector;
  --gpib_edm1_clock_2_in_end_xfer assignment, which is an e_assign
  gpib_edm1_clock_2_in_end_xfer <= NOT ((gpib_edm1_clock_2_in_waits_for_read OR gpib_edm1_clock_2_in_waits_for_write));
  --end_xfer_arb_share_counter_term_gpib_edm1_clock_2_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gpib_edm1_clock_2_in <= gpib_edm1_clock_2_in_end_xfer AND (((NOT gpib_edm1_clock_2_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gpib_edm1_clock_2_in_arb_share_counter arbitration counter enable, which is an e_assign
  gpib_edm1_clock_2_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gpib_edm1_clock_2_in AND gpib_edm1_clock_2_in_allgrants)) OR ((end_xfer_arb_share_counter_term_gpib_edm1_clock_2_in AND NOT gpib_edm1_clock_2_in_non_bursting_master_requests));
  --gpib_edm1_clock_2_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_2_in_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gpib_edm1_clock_2_in_arb_counter_enable) = '1' then 
        gpib_edm1_clock_2_in_arb_share_counter <= gpib_edm1_clock_2_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_2_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_2_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gpib_edm1_clock_2_in_master_qreq_vector AND end_xfer_arb_share_counter_term_gpib_edm1_clock_2_in)) OR ((end_xfer_arb_share_counter_term_gpib_edm1_clock_2_in AND NOT gpib_edm1_clock_2_in_non_bursting_master_requests)))) = '1' then 
        gpib_edm1_clock_2_in_slavearbiterlockenable <= gpib_edm1_clock_2_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 gpib_edm1_clock_2/in arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= gpib_edm1_clock_2_in_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --gpib_edm1_clock_2_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gpib_edm1_clock_2_in_slavearbiterlockenable2 <= gpib_edm1_clock_2_in_arb_share_counter_next_value;
  --clock_crossing_0/m1 gpib_edm1_clock_2/in arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= gpib_edm1_clock_2_in_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --gpib_edm1_clock_2_in_any_continuerequest at least one master continues requesting, which is an e_assign
  gpib_edm1_clock_2_in_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in <= internal_clock_crossing_0_m1_requests_gpib_edm1_clock_2_in AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in, which is an e_mux
  clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in <= (internal_clock_crossing_0_m1_granted_gpib_edm1_clock_2_in AND clock_crossing_0_m1_read) AND NOT gpib_edm1_clock_2_in_waits_for_read;
  --gpib_edm1_clock_2_in_writedata mux, which is an e_mux
  gpib_edm1_clock_2_in_writedata <= clock_crossing_0_m1_writedata (15 DOWNTO 0);
  --assign gpib_edm1_clock_2_in_endofpacket_from_sa = gpib_edm1_clock_2_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpib_edm1_clock_2_in_endofpacket_from_sa <= gpib_edm1_clock_2_in_endofpacket;
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_gpib_edm1_clock_2_in <= internal_clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in;
  --clock_crossing_0/m1 saved-grant gpib_edm1_clock_2/in, which is an e_assign
  clock_crossing_0_m1_saved_grant_gpib_edm1_clock_2_in <= internal_clock_crossing_0_m1_requests_gpib_edm1_clock_2_in;
  --allow new arb cycle for gpib_edm1_clock_2/in, which is an e_assign
  gpib_edm1_clock_2_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gpib_edm1_clock_2_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gpib_edm1_clock_2_in_master_qreq_vector <= std_logic'('1');
  --gpib_edm1_clock_2_in_reset_n assignment, which is an e_assign
  gpib_edm1_clock_2_in_reset_n <= reset_n;
  --gpib_edm1_clock_2_in_firsttransfer first transaction, which is an e_assign
  gpib_edm1_clock_2_in_firsttransfer <= A_WE_StdLogic((std_logic'(gpib_edm1_clock_2_in_begins_xfer) = '1'), gpib_edm1_clock_2_in_unreg_firsttransfer, gpib_edm1_clock_2_in_reg_firsttransfer);
  --gpib_edm1_clock_2_in_unreg_firsttransfer first transaction, which is an e_assign
  gpib_edm1_clock_2_in_unreg_firsttransfer <= NOT ((gpib_edm1_clock_2_in_slavearbiterlockenable AND gpib_edm1_clock_2_in_any_continuerequest));
  --gpib_edm1_clock_2_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_2_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gpib_edm1_clock_2_in_begins_xfer) = '1' then 
        gpib_edm1_clock_2_in_reg_firsttransfer <= gpib_edm1_clock_2_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_2_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gpib_edm1_clock_2_in_beginbursttransfer_internal <= gpib_edm1_clock_2_in_begins_xfer;
  --gpib_edm1_clock_2_in_read assignment, which is an e_mux
  gpib_edm1_clock_2_in_read <= internal_clock_crossing_0_m1_granted_gpib_edm1_clock_2_in AND clock_crossing_0_m1_read;
  --gpib_edm1_clock_2_in_write assignment, which is an e_mux
  gpib_edm1_clock_2_in_write <= internal_clock_crossing_0_m1_granted_gpib_edm1_clock_2_in AND clock_crossing_0_m1_write;
  --gpib_edm1_clock_2_in_address mux, which is an e_mux
  gpib_edm1_clock_2_in_address <= clock_crossing_0_m1_address_to_slave (3 DOWNTO 0);
  --slaveid gpib_edm1_clock_2_in_nativeaddress nativeaddress mux, which is an e_mux
  gpib_edm1_clock_2_in_nativeaddress <= clock_crossing_0_m1_nativeaddress (2 DOWNTO 0);
  --d1_gpib_edm1_clock_2_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gpib_edm1_clock_2_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gpib_edm1_clock_2_in_end_xfer <= gpib_edm1_clock_2_in_end_xfer;
    end if;

  end process;

  --gpib_edm1_clock_2_in_waits_for_read in a cycle, which is an e_mux
  gpib_edm1_clock_2_in_waits_for_read <= gpib_edm1_clock_2_in_in_a_read_cycle AND internal_gpib_edm1_clock_2_in_waitrequest_from_sa;
  --gpib_edm1_clock_2_in_in_a_read_cycle assignment, which is an e_assign
  gpib_edm1_clock_2_in_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_gpib_edm1_clock_2_in AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gpib_edm1_clock_2_in_in_a_read_cycle;
  --gpib_edm1_clock_2_in_waits_for_write in a cycle, which is an e_mux
  gpib_edm1_clock_2_in_waits_for_write <= gpib_edm1_clock_2_in_in_a_write_cycle AND internal_gpib_edm1_clock_2_in_waitrequest_from_sa;
  --gpib_edm1_clock_2_in_in_a_write_cycle assignment, which is an e_assign
  gpib_edm1_clock_2_in_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_gpib_edm1_clock_2_in AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gpib_edm1_clock_2_in_in_a_write_cycle;
  wait_for_gpib_edm1_clock_2_in_counter <= std_logic'('0');
  --gpib_edm1_clock_2_in_byteenable byte enable port mux, which is an e_mux
  gpib_edm1_clock_2_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_clock_crossing_0_m1_granted_gpib_edm1_clock_2_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (clock_crossing_0_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_gpib_edm1_clock_2_in <= internal_clock_crossing_0_m1_granted_gpib_edm1_clock_2_in;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in <= internal_clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_gpib_edm1_clock_2_in <= internal_clock_crossing_0_m1_requests_gpib_edm1_clock_2_in;
  --vhdl renameroo for output signals
  gpib_edm1_clock_2_in_waitrequest_from_sa <= internal_gpib_edm1_clock_2_in_waitrequest_from_sa;
--synthesis translate_off
    --gpib_edm1_clock_2/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity gpib_edm1_clock_2_out_arbitrator is 
        port (
              -- inputs:
                 signal ad7928_spi_control_port_endofpacket_from_sa : IN STD_LOGIC;
                 signal ad7928_spi_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_ad7928_spi_control_port_end_xfer : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_2_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gpib_edm1_clock_2_out_granted_ad7928_spi_control_port : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_out_read : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_out_read_data_valid_ad7928_spi_control_port : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_out_requests_ad7928_spi_control_port : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_out_write : IN STD_LOGIC;
                 signal gpib_edm1_clock_2_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal gpib_edm1_clock_2_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_2_out_endofpacket : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_2_out_reset_n : OUT STD_LOGIC;
                 signal gpib_edm1_clock_2_out_waitrequest : OUT STD_LOGIC
              );
end entity gpib_edm1_clock_2_out_arbitrator;


architecture europa of gpib_edm1_clock_2_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_2_out_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_edm1_clock_2_out_read_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_run :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_write_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_gpib_edm1_clock_2_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_gpib_edm1_clock_2_out_waitrequest :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port OR NOT ((gpib_edm1_clock_2_out_read OR gpib_edm1_clock_2_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_ad7928_spi_control_port_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((gpib_edm1_clock_2_out_read OR gpib_edm1_clock_2_out_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port OR NOT ((gpib_edm1_clock_2_out_read OR gpib_edm1_clock_2_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_ad7928_spi_control_port_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((gpib_edm1_clock_2_out_read OR gpib_edm1_clock_2_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  gpib_edm1_clock_2_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_gpib_edm1_clock_2_out_address_to_slave <= gpib_edm1_clock_2_out_address;
  --gpib_edm1_clock_2/out readdata mux, which is an e_mux
  gpib_edm1_clock_2_out_readdata <= ad7928_spi_control_port_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_gpib_edm1_clock_2_out_waitrequest <= NOT gpib_edm1_clock_2_out_run;
  --gpib_edm1_clock_2_out_reset_n assignment, which is an e_assign
  gpib_edm1_clock_2_out_reset_n <= reset_n;
  --mux gpib_edm1_clock_2_out_endofpacket, which is an e_mux
  gpib_edm1_clock_2_out_endofpacket <= ad7928_spi_control_port_endofpacket_from_sa;
  --vhdl renameroo for output signals
  gpib_edm1_clock_2_out_address_to_slave <= internal_gpib_edm1_clock_2_out_address_to_slave;
  --vhdl renameroo for output signals
  gpib_edm1_clock_2_out_waitrequest <= internal_gpib_edm1_clock_2_out_waitrequest;
--synthesis translate_off
    --gpib_edm1_clock_2_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_2_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_2_out_address_last_time <= gpib_edm1_clock_2_out_address;
      end if;

    end process;

    --gpib_edm1_clock_2/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_gpib_edm1_clock_2_out_waitrequest AND ((gpib_edm1_clock_2_out_read OR gpib_edm1_clock_2_out_write));
      end if;

    end process;

    --gpib_edm1_clock_2_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line40 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_2_out_address /= gpib_edm1_clock_2_out_address_last_time))))) = '1' then 
          write(write_line40, now);
          write(write_line40, string'(": "));
          write(write_line40, string'("gpib_edm1_clock_2_out_address did not heed wait!!!"));
          write(output, write_line40.all);
          deallocate (write_line40);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_2_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_2_out_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_2_out_byteenable_last_time <= gpib_edm1_clock_2_out_byteenable;
      end if;

    end process;

    --gpib_edm1_clock_2_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line41 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_2_out_byteenable /= gpib_edm1_clock_2_out_byteenable_last_time))))) = '1' then 
          write(write_line41, now);
          write(write_line41, string'(": "));
          write(write_line41, string'("gpib_edm1_clock_2_out_byteenable did not heed wait!!!"));
          write(output, write_line41.all);
          deallocate (write_line41);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_2_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_2_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_2_out_read_last_time <= gpib_edm1_clock_2_out_read;
      end if;

    end process;

    --gpib_edm1_clock_2_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line42 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(gpib_edm1_clock_2_out_read) /= std_logic'(gpib_edm1_clock_2_out_read_last_time)))))) = '1' then 
          write(write_line42, now);
          write(write_line42, string'(": "));
          write(write_line42, string'("gpib_edm1_clock_2_out_read did not heed wait!!!"));
          write(output, write_line42.all);
          deallocate (write_line42);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_2_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_2_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_2_out_write_last_time <= gpib_edm1_clock_2_out_write;
      end if;

    end process;

    --gpib_edm1_clock_2_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line43 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(gpib_edm1_clock_2_out_write) /= std_logic'(gpib_edm1_clock_2_out_write_last_time)))))) = '1' then 
          write(write_line43, now);
          write(write_line43, string'(": "));
          write(write_line43, string'("gpib_edm1_clock_2_out_write did not heed wait!!!"));
          write(output, write_line43.all);
          deallocate (write_line43);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_2_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_2_out_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_2_out_writedata_last_time <= gpib_edm1_clock_2_out_writedata;
      end if;

    end process;

    --gpib_edm1_clock_2_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line44 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_2_out_writedata /= gpib_edm1_clock_2_out_writedata_last_time)))) AND gpib_edm1_clock_2_out_write)) = '1' then 
          write(write_line44, now);
          write(write_line44, string'(": "));
          write(write_line44, string'("gpib_edm1_clock_2_out_writedata did not heed wait!!!"));
          write(output, write_line44.all);
          deallocate (write_line44);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_edm1_clock_3_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpib_edm1_clock_3_in_endofpacket : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_3_in_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_m1_granted_gpib_edm1_clock_3_in : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_gpib_edm1_clock_3_in : OUT STD_LOGIC;
                 signal d1_gpib_edm1_clock_3_in_end_xfer : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_3_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gpib_edm1_clock_3_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal gpib_edm1_clock_3_in_read : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_3_in_reset_n : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_in_write : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity gpib_edm1_clock_3_in_arbitrator;


architecture europa of gpib_edm1_clock_3_in_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_gpib_edm1_clock_3_in :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gpib_edm1_clock_3_in :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_allgrants :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_allow_new_arb_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_any_continuerequest :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_arb_counter_enable :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_arb_share_counter :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_arb_share_counter_next_value :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_arb_share_set_values :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_beginbursttransfer_internal :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_begins_xfer :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_end_xfer :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_grant_vector :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_in_a_read_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_in_a_write_cycle :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_master_qreq_vector :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_non_bursting_master_requests :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_reg_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_slavearbiterlockenable :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_unreg_firsttransfer :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_waits_for_read :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_gpib_edm1_clock_3_in :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_gpib_edm1_clock_3_in :  STD_LOGIC;
                signal internal_gpib_edm1_clock_3_in_waitrequest_from_sa :  STD_LOGIC;
                signal wait_for_gpib_edm1_clock_3_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gpib_edm1_clock_3_in_end_xfer;
    end if;

  end process;

  gpib_edm1_clock_3_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in);
  --assign gpib_edm1_clock_3_in_readdata_from_sa = gpib_edm1_clock_3_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpib_edm1_clock_3_in_readdata_from_sa <= gpib_edm1_clock_3_in_readdata;
  internal_clock_crossing_0_m1_requests_gpib_edm1_clock_3_in <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(7 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("10000000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --assign gpib_edm1_clock_3_in_waitrequest_from_sa = gpib_edm1_clock_3_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_gpib_edm1_clock_3_in_waitrequest_from_sa <= gpib_edm1_clock_3_in_waitrequest;
  --gpib_edm1_clock_3_in_arb_share_counter set values, which is an e_mux
  gpib_edm1_clock_3_in_arb_share_set_values <= std_logic'('1');
  --gpib_edm1_clock_3_in_non_bursting_master_requests mux, which is an e_mux
  gpib_edm1_clock_3_in_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_gpib_edm1_clock_3_in;
  --gpib_edm1_clock_3_in_any_bursting_master_saved_grant mux, which is an e_mux
  gpib_edm1_clock_3_in_any_bursting_master_saved_grant <= std_logic'('0');
  --gpib_edm1_clock_3_in_arb_share_counter_next_value assignment, which is an e_assign
  gpib_edm1_clock_3_in_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gpib_edm1_clock_3_in_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_edm1_clock_3_in_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gpib_edm1_clock_3_in_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_edm1_clock_3_in_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gpib_edm1_clock_3_in_allgrants all slave grants, which is an e_mux
  gpib_edm1_clock_3_in_allgrants <= gpib_edm1_clock_3_in_grant_vector;
  --gpib_edm1_clock_3_in_end_xfer assignment, which is an e_assign
  gpib_edm1_clock_3_in_end_xfer <= NOT ((gpib_edm1_clock_3_in_waits_for_read OR gpib_edm1_clock_3_in_waits_for_write));
  --end_xfer_arb_share_counter_term_gpib_edm1_clock_3_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gpib_edm1_clock_3_in <= gpib_edm1_clock_3_in_end_xfer AND (((NOT gpib_edm1_clock_3_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gpib_edm1_clock_3_in_arb_share_counter arbitration counter enable, which is an e_assign
  gpib_edm1_clock_3_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gpib_edm1_clock_3_in AND gpib_edm1_clock_3_in_allgrants)) OR ((end_xfer_arb_share_counter_term_gpib_edm1_clock_3_in AND NOT gpib_edm1_clock_3_in_non_bursting_master_requests));
  --gpib_edm1_clock_3_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_3_in_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gpib_edm1_clock_3_in_arb_counter_enable) = '1' then 
        gpib_edm1_clock_3_in_arb_share_counter <= gpib_edm1_clock_3_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_3_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_3_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gpib_edm1_clock_3_in_master_qreq_vector AND end_xfer_arb_share_counter_term_gpib_edm1_clock_3_in)) OR ((end_xfer_arb_share_counter_term_gpib_edm1_clock_3_in AND NOT gpib_edm1_clock_3_in_non_bursting_master_requests)))) = '1' then 
        gpib_edm1_clock_3_in_slavearbiterlockenable <= gpib_edm1_clock_3_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 gpib_edm1_clock_3/in arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= gpib_edm1_clock_3_in_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --gpib_edm1_clock_3_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gpib_edm1_clock_3_in_slavearbiterlockenable2 <= gpib_edm1_clock_3_in_arb_share_counter_next_value;
  --clock_crossing_0/m1 gpib_edm1_clock_3/in arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= gpib_edm1_clock_3_in_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --gpib_edm1_clock_3_in_any_continuerequest at least one master continues requesting, which is an e_assign
  gpib_edm1_clock_3_in_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in <= internal_clock_crossing_0_m1_requests_gpib_edm1_clock_3_in AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in, which is an e_mux
  clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in <= (internal_clock_crossing_0_m1_granted_gpib_edm1_clock_3_in AND clock_crossing_0_m1_read) AND NOT gpib_edm1_clock_3_in_waits_for_read;
  --gpib_edm1_clock_3_in_writedata mux, which is an e_mux
  gpib_edm1_clock_3_in_writedata <= clock_crossing_0_m1_writedata (15 DOWNTO 0);
  --assign gpib_edm1_clock_3_in_endofpacket_from_sa = gpib_edm1_clock_3_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpib_edm1_clock_3_in_endofpacket_from_sa <= gpib_edm1_clock_3_in_endofpacket;
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_gpib_edm1_clock_3_in <= internal_clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in;
  --clock_crossing_0/m1 saved-grant gpib_edm1_clock_3/in, which is an e_assign
  clock_crossing_0_m1_saved_grant_gpib_edm1_clock_3_in <= internal_clock_crossing_0_m1_requests_gpib_edm1_clock_3_in;
  --allow new arb cycle for gpib_edm1_clock_3/in, which is an e_assign
  gpib_edm1_clock_3_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gpib_edm1_clock_3_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gpib_edm1_clock_3_in_master_qreq_vector <= std_logic'('1');
  --gpib_edm1_clock_3_in_reset_n assignment, which is an e_assign
  gpib_edm1_clock_3_in_reset_n <= reset_n;
  --gpib_edm1_clock_3_in_firsttransfer first transaction, which is an e_assign
  gpib_edm1_clock_3_in_firsttransfer <= A_WE_StdLogic((std_logic'(gpib_edm1_clock_3_in_begins_xfer) = '1'), gpib_edm1_clock_3_in_unreg_firsttransfer, gpib_edm1_clock_3_in_reg_firsttransfer);
  --gpib_edm1_clock_3_in_unreg_firsttransfer first transaction, which is an e_assign
  gpib_edm1_clock_3_in_unreg_firsttransfer <= NOT ((gpib_edm1_clock_3_in_slavearbiterlockenable AND gpib_edm1_clock_3_in_any_continuerequest));
  --gpib_edm1_clock_3_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_3_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gpib_edm1_clock_3_in_begins_xfer) = '1' then 
        gpib_edm1_clock_3_in_reg_firsttransfer <= gpib_edm1_clock_3_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_3_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gpib_edm1_clock_3_in_beginbursttransfer_internal <= gpib_edm1_clock_3_in_begins_xfer;
  --gpib_edm1_clock_3_in_read assignment, which is an e_mux
  gpib_edm1_clock_3_in_read <= internal_clock_crossing_0_m1_granted_gpib_edm1_clock_3_in AND clock_crossing_0_m1_read;
  --gpib_edm1_clock_3_in_write assignment, which is an e_mux
  gpib_edm1_clock_3_in_write <= internal_clock_crossing_0_m1_granted_gpib_edm1_clock_3_in AND clock_crossing_0_m1_write;
  --gpib_edm1_clock_3_in_address mux, which is an e_mux
  gpib_edm1_clock_3_in_address <= clock_crossing_0_m1_address_to_slave (3 DOWNTO 0);
  --slaveid gpib_edm1_clock_3_in_nativeaddress nativeaddress mux, which is an e_mux
  gpib_edm1_clock_3_in_nativeaddress <= clock_crossing_0_m1_nativeaddress (2 DOWNTO 0);
  --d1_gpib_edm1_clock_3_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gpib_edm1_clock_3_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gpib_edm1_clock_3_in_end_xfer <= gpib_edm1_clock_3_in_end_xfer;
    end if;

  end process;

  --gpib_edm1_clock_3_in_waits_for_read in a cycle, which is an e_mux
  gpib_edm1_clock_3_in_waits_for_read <= gpib_edm1_clock_3_in_in_a_read_cycle AND internal_gpib_edm1_clock_3_in_waitrequest_from_sa;
  --gpib_edm1_clock_3_in_in_a_read_cycle assignment, which is an e_assign
  gpib_edm1_clock_3_in_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_gpib_edm1_clock_3_in AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gpib_edm1_clock_3_in_in_a_read_cycle;
  --gpib_edm1_clock_3_in_waits_for_write in a cycle, which is an e_mux
  gpib_edm1_clock_3_in_waits_for_write <= gpib_edm1_clock_3_in_in_a_write_cycle AND internal_gpib_edm1_clock_3_in_waitrequest_from_sa;
  --gpib_edm1_clock_3_in_in_a_write_cycle assignment, which is an e_assign
  gpib_edm1_clock_3_in_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_gpib_edm1_clock_3_in AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gpib_edm1_clock_3_in_in_a_write_cycle;
  wait_for_gpib_edm1_clock_3_in_counter <= std_logic'('0');
  --gpib_edm1_clock_3_in_byteenable byte enable port mux, which is an e_mux
  gpib_edm1_clock_3_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_clock_crossing_0_m1_granted_gpib_edm1_clock_3_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (clock_crossing_0_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_gpib_edm1_clock_3_in <= internal_clock_crossing_0_m1_granted_gpib_edm1_clock_3_in;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in <= internal_clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_gpib_edm1_clock_3_in <= internal_clock_crossing_0_m1_requests_gpib_edm1_clock_3_in;
  --vhdl renameroo for output signals
  gpib_edm1_clock_3_in_waitrequest_from_sa <= internal_gpib_edm1_clock_3_in_waitrequest_from_sa;
--synthesis translate_off
    --gpib_edm1_clock_3/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity gpib_edm1_clock_3_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_dac_ad5308_spi_control_port_end_xfer : IN STD_LOGIC;
                 signal dac_ad5308_spi_control_port_endofpacket_from_sa : IN STD_LOGIC;
                 signal dac_ad5308_spi_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_3_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_3_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_out_read : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_out_read_data_valid_dac_ad5308_spi_control_port : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_out_write : IN STD_LOGIC;
                 signal gpib_edm1_clock_3_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal gpib_edm1_clock_3_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_3_out_endofpacket : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal gpib_edm1_clock_3_out_reset_n : OUT STD_LOGIC;
                 signal gpib_edm1_clock_3_out_waitrequest : OUT STD_LOGIC
              );
end entity gpib_edm1_clock_3_out_arbitrator;


architecture europa of gpib_edm1_clock_3_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_3_out_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_edm1_clock_3_out_read_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_run :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_write_last_time :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_gpib_edm1_clock_3_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_gpib_edm1_clock_3_out_waitrequest :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port OR NOT ((gpib_edm1_clock_3_out_read OR gpib_edm1_clock_3_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_dac_ad5308_spi_control_port_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((gpib_edm1_clock_3_out_read OR gpib_edm1_clock_3_out_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port OR NOT ((gpib_edm1_clock_3_out_read OR gpib_edm1_clock_3_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_dac_ad5308_spi_control_port_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((gpib_edm1_clock_3_out_read OR gpib_edm1_clock_3_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  gpib_edm1_clock_3_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_gpib_edm1_clock_3_out_address_to_slave <= gpib_edm1_clock_3_out_address;
  --gpib_edm1_clock_3/out readdata mux, which is an e_mux
  gpib_edm1_clock_3_out_readdata <= dac_ad5308_spi_control_port_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_gpib_edm1_clock_3_out_waitrequest <= NOT gpib_edm1_clock_3_out_run;
  --gpib_edm1_clock_3_out_reset_n assignment, which is an e_assign
  gpib_edm1_clock_3_out_reset_n <= reset_n;
  --mux gpib_edm1_clock_3_out_endofpacket, which is an e_mux
  gpib_edm1_clock_3_out_endofpacket <= dac_ad5308_spi_control_port_endofpacket_from_sa;
  --vhdl renameroo for output signals
  gpib_edm1_clock_3_out_address_to_slave <= internal_gpib_edm1_clock_3_out_address_to_slave;
  --vhdl renameroo for output signals
  gpib_edm1_clock_3_out_waitrequest <= internal_gpib_edm1_clock_3_out_waitrequest;
--synthesis translate_off
    --gpib_edm1_clock_3_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_3_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_3_out_address_last_time <= gpib_edm1_clock_3_out_address;
      end if;

    end process;

    --gpib_edm1_clock_3/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_gpib_edm1_clock_3_out_waitrequest AND ((gpib_edm1_clock_3_out_read OR gpib_edm1_clock_3_out_write));
      end if;

    end process;

    --gpib_edm1_clock_3_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line45 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_3_out_address /= gpib_edm1_clock_3_out_address_last_time))))) = '1' then 
          write(write_line45, now);
          write(write_line45, string'(": "));
          write(write_line45, string'("gpib_edm1_clock_3_out_address did not heed wait!!!"));
          write(output, write_line45.all);
          deallocate (write_line45);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_3_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_3_out_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_3_out_byteenable_last_time <= gpib_edm1_clock_3_out_byteenable;
      end if;

    end process;

    --gpib_edm1_clock_3_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line46 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_3_out_byteenable /= gpib_edm1_clock_3_out_byteenable_last_time))))) = '1' then 
          write(write_line46, now);
          write(write_line46, string'(": "));
          write(write_line46, string'("gpib_edm1_clock_3_out_byteenable did not heed wait!!!"));
          write(output, write_line46.all);
          deallocate (write_line46);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_3_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_3_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_3_out_read_last_time <= gpib_edm1_clock_3_out_read;
      end if;

    end process;

    --gpib_edm1_clock_3_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line47 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(gpib_edm1_clock_3_out_read) /= std_logic'(gpib_edm1_clock_3_out_read_last_time)))))) = '1' then 
          write(write_line47, now);
          write(write_line47, string'(": "));
          write(write_line47, string'("gpib_edm1_clock_3_out_read did not heed wait!!!"));
          write(output, write_line47.all);
          deallocate (write_line47);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_3_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_3_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_3_out_write_last_time <= gpib_edm1_clock_3_out_write;
      end if;

    end process;

    --gpib_edm1_clock_3_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line48 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(gpib_edm1_clock_3_out_write) /= std_logic'(gpib_edm1_clock_3_out_write_last_time)))))) = '1' then 
          write(write_line48, now);
          write(write_line48, string'(": "));
          write(write_line48, string'("gpib_edm1_clock_3_out_write did not heed wait!!!"));
          write(output, write_line48.all);
          deallocate (write_line48);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --gpib_edm1_clock_3_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        gpib_edm1_clock_3_out_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        gpib_edm1_clock_3_out_writedata_last_time <= gpib_edm1_clock_3_out_writedata;
      end if;

    end process;

    --gpib_edm1_clock_3_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line49 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((gpib_edm1_clock_3_out_writedata /= gpib_edm1_clock_3_out_writedata_last_time)))) AND gpib_edm1_clock_3_out_write)) = '1' then 
          write(write_line49, now);
          write(write_line49, string'(": "));
          write(write_line49, string'("gpib_edm1_clock_3_out_writedata did not heed wait!!!"));
          write(output, write_line49.all);
          deallocate (write_line49);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_leds_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpib_leds_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_m1_granted_gpib_leds_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_gpib_leds_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_gpib_leds_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_gpib_leds_s1 : OUT STD_LOGIC;
                 signal d1_gpib_leds_s1_end_xfer : OUT STD_LOGIC;
                 signal gpib_leds_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gpib_leds_s1_chipselect : OUT STD_LOGIC;
                 signal gpib_leds_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gpib_leds_s1_reset_n : OUT STD_LOGIC;
                 signal gpib_leds_s1_write_n : OUT STD_LOGIC;
                 signal gpib_leds_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity gpib_leds_s1_arbitrator;


architecture europa of gpib_leds_s1_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_gpib_leds_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gpib_leds_s1 :  STD_LOGIC;
                signal gpib_leds_s1_allgrants :  STD_LOGIC;
                signal gpib_leds_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal gpib_leds_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gpib_leds_s1_any_continuerequest :  STD_LOGIC;
                signal gpib_leds_s1_arb_counter_enable :  STD_LOGIC;
                signal gpib_leds_s1_arb_share_counter :  STD_LOGIC;
                signal gpib_leds_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal gpib_leds_s1_arb_share_set_values :  STD_LOGIC;
                signal gpib_leds_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal gpib_leds_s1_begins_xfer :  STD_LOGIC;
                signal gpib_leds_s1_end_xfer :  STD_LOGIC;
                signal gpib_leds_s1_firsttransfer :  STD_LOGIC;
                signal gpib_leds_s1_grant_vector :  STD_LOGIC;
                signal gpib_leds_s1_in_a_read_cycle :  STD_LOGIC;
                signal gpib_leds_s1_in_a_write_cycle :  STD_LOGIC;
                signal gpib_leds_s1_master_qreq_vector :  STD_LOGIC;
                signal gpib_leds_s1_non_bursting_master_requests :  STD_LOGIC;
                signal gpib_leds_s1_pretend_byte_enable :  STD_LOGIC;
                signal gpib_leds_s1_reg_firsttransfer :  STD_LOGIC;
                signal gpib_leds_s1_slavearbiterlockenable :  STD_LOGIC;
                signal gpib_leds_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal gpib_leds_s1_unreg_firsttransfer :  STD_LOGIC;
                signal gpib_leds_s1_waits_for_read :  STD_LOGIC;
                signal gpib_leds_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_gpib_leds_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_gpib_leds_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_gpib_leds_s1 :  STD_LOGIC;
                signal wait_for_gpib_leds_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gpib_leds_s1_end_xfer;
    end if;

  end process;

  gpib_leds_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_gpib_leds_s1);
  --assign gpib_leds_s1_readdata_from_sa = gpib_leds_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpib_leds_s1_readdata_from_sa <= gpib_leds_s1_readdata;
  internal_clock_crossing_0_m1_requests_gpib_leds_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(7 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10110000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --gpib_leds_s1_arb_share_counter set values, which is an e_mux
  gpib_leds_s1_arb_share_set_values <= std_logic'('1');
  --gpib_leds_s1_non_bursting_master_requests mux, which is an e_mux
  gpib_leds_s1_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_gpib_leds_s1;
  --gpib_leds_s1_any_bursting_master_saved_grant mux, which is an e_mux
  gpib_leds_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --gpib_leds_s1_arb_share_counter_next_value assignment, which is an e_assign
  gpib_leds_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gpib_leds_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_leds_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gpib_leds_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_leds_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gpib_leds_s1_allgrants all slave grants, which is an e_mux
  gpib_leds_s1_allgrants <= gpib_leds_s1_grant_vector;
  --gpib_leds_s1_end_xfer assignment, which is an e_assign
  gpib_leds_s1_end_xfer <= NOT ((gpib_leds_s1_waits_for_read OR gpib_leds_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_gpib_leds_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gpib_leds_s1 <= gpib_leds_s1_end_xfer AND (((NOT gpib_leds_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gpib_leds_s1_arb_share_counter arbitration counter enable, which is an e_assign
  gpib_leds_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gpib_leds_s1 AND gpib_leds_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_gpib_leds_s1 AND NOT gpib_leds_s1_non_bursting_master_requests));
  --gpib_leds_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_leds_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gpib_leds_s1_arb_counter_enable) = '1' then 
        gpib_leds_s1_arb_share_counter <= gpib_leds_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpib_leds_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_leds_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gpib_leds_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_gpib_leds_s1)) OR ((end_xfer_arb_share_counter_term_gpib_leds_s1 AND NOT gpib_leds_s1_non_bursting_master_requests)))) = '1' then 
        gpib_leds_s1_slavearbiterlockenable <= gpib_leds_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 gpib_leds/s1 arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= gpib_leds_s1_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --gpib_leds_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gpib_leds_s1_slavearbiterlockenable2 <= gpib_leds_s1_arb_share_counter_next_value;
  --clock_crossing_0/m1 gpib_leds/s1 arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= gpib_leds_s1_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --gpib_leds_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  gpib_leds_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_gpib_leds_s1 <= internal_clock_crossing_0_m1_requests_gpib_leds_s1 AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_gpib_leds_s1, which is an e_mux
  clock_crossing_0_m1_read_data_valid_gpib_leds_s1 <= (internal_clock_crossing_0_m1_granted_gpib_leds_s1 AND clock_crossing_0_m1_read) AND NOT gpib_leds_s1_waits_for_read;
  --gpib_leds_s1_writedata mux, which is an e_mux
  gpib_leds_s1_writedata <= clock_crossing_0_m1_writedata (7 DOWNTO 0);
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_gpib_leds_s1 <= internal_clock_crossing_0_m1_qualified_request_gpib_leds_s1;
  --clock_crossing_0/m1 saved-grant gpib_leds/s1, which is an e_assign
  clock_crossing_0_m1_saved_grant_gpib_leds_s1 <= internal_clock_crossing_0_m1_requests_gpib_leds_s1;
  --allow new arb cycle for gpib_leds/s1, which is an e_assign
  gpib_leds_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gpib_leds_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gpib_leds_s1_master_qreq_vector <= std_logic'('1');
  --gpib_leds_s1_reset_n assignment, which is an e_assign
  gpib_leds_s1_reset_n <= reset_n;
  gpib_leds_s1_chipselect <= internal_clock_crossing_0_m1_granted_gpib_leds_s1;
  --gpib_leds_s1_firsttransfer first transaction, which is an e_assign
  gpib_leds_s1_firsttransfer <= A_WE_StdLogic((std_logic'(gpib_leds_s1_begins_xfer) = '1'), gpib_leds_s1_unreg_firsttransfer, gpib_leds_s1_reg_firsttransfer);
  --gpib_leds_s1_unreg_firsttransfer first transaction, which is an e_assign
  gpib_leds_s1_unreg_firsttransfer <= NOT ((gpib_leds_s1_slavearbiterlockenable AND gpib_leds_s1_any_continuerequest));
  --gpib_leds_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_leds_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gpib_leds_s1_begins_xfer) = '1' then 
        gpib_leds_s1_reg_firsttransfer <= gpib_leds_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gpib_leds_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gpib_leds_s1_beginbursttransfer_internal <= gpib_leds_s1_begins_xfer;
  --~gpib_leds_s1_write_n assignment, which is an e_mux
  gpib_leds_s1_write_n <= NOT ((((internal_clock_crossing_0_m1_granted_gpib_leds_s1 AND clock_crossing_0_m1_write)) AND gpib_leds_s1_pretend_byte_enable));
  --gpib_leds_s1_address mux, which is an e_mux
  gpib_leds_s1_address <= clock_crossing_0_m1_nativeaddress (1 DOWNTO 0);
  --d1_gpib_leds_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gpib_leds_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gpib_leds_s1_end_xfer <= gpib_leds_s1_end_xfer;
    end if;

  end process;

  --gpib_leds_s1_waits_for_read in a cycle, which is an e_mux
  gpib_leds_s1_waits_for_read <= gpib_leds_s1_in_a_read_cycle AND gpib_leds_s1_begins_xfer;
  --gpib_leds_s1_in_a_read_cycle assignment, which is an e_assign
  gpib_leds_s1_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_gpib_leds_s1 AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gpib_leds_s1_in_a_read_cycle;
  --gpib_leds_s1_waits_for_write in a cycle, which is an e_mux
  gpib_leds_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpib_leds_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --gpib_leds_s1_in_a_write_cycle assignment, which is an e_assign
  gpib_leds_s1_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_gpib_leds_s1 AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gpib_leds_s1_in_a_write_cycle;
  wait_for_gpib_leds_s1_counter <= std_logic'('0');
  --gpib_leds_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  gpib_leds_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_clock_crossing_0_m1_granted_gpib_leds_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (clock_crossing_0_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_gpib_leds_s1 <= internal_clock_crossing_0_m1_granted_gpib_leds_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_gpib_leds_s1 <= internal_clock_crossing_0_m1_qualified_request_gpib_leds_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_gpib_leds_s1 <= internal_clock_crossing_0_m1_requests_gpib_leds_s1;
--synthesis translate_off
    --gpib_leds/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpio1_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpio1_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_m1_granted_gpio1_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_gpio1_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_gpio1_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_gpio1_s1 : OUT STD_LOGIC;
                 signal d1_gpio1_s1_end_xfer : OUT STD_LOGIC;
                 signal gpio1_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal gpio1_s1_chipselect : OUT STD_LOGIC;
                 signal gpio1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gpio1_s1_reset_n : OUT STD_LOGIC;
                 signal gpio1_s1_write_n : OUT STD_LOGIC;
                 signal gpio1_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity gpio1_s1_arbitrator;


architecture europa of gpio1_s1_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_gpio1_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gpio1_s1 :  STD_LOGIC;
                signal gpio1_s1_allgrants :  STD_LOGIC;
                signal gpio1_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal gpio1_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gpio1_s1_any_continuerequest :  STD_LOGIC;
                signal gpio1_s1_arb_counter_enable :  STD_LOGIC;
                signal gpio1_s1_arb_share_counter :  STD_LOGIC;
                signal gpio1_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal gpio1_s1_arb_share_set_values :  STD_LOGIC;
                signal gpio1_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal gpio1_s1_begins_xfer :  STD_LOGIC;
                signal gpio1_s1_end_xfer :  STD_LOGIC;
                signal gpio1_s1_firsttransfer :  STD_LOGIC;
                signal gpio1_s1_grant_vector :  STD_LOGIC;
                signal gpio1_s1_in_a_read_cycle :  STD_LOGIC;
                signal gpio1_s1_in_a_write_cycle :  STD_LOGIC;
                signal gpio1_s1_master_qreq_vector :  STD_LOGIC;
                signal gpio1_s1_non_bursting_master_requests :  STD_LOGIC;
                signal gpio1_s1_pretend_byte_enable :  STD_LOGIC;
                signal gpio1_s1_reg_firsttransfer :  STD_LOGIC;
                signal gpio1_s1_slavearbiterlockenable :  STD_LOGIC;
                signal gpio1_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal gpio1_s1_unreg_firsttransfer :  STD_LOGIC;
                signal gpio1_s1_waits_for_read :  STD_LOGIC;
                signal gpio1_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_gpio1_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_gpio1_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_gpio1_s1 :  STD_LOGIC;
                signal wait_for_gpio1_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gpio1_s1_end_xfer;
    end if;

  end process;

  gpio1_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_gpio1_s1);
  --assign gpio1_s1_readdata_from_sa = gpio1_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpio1_s1_readdata_from_sa <= gpio1_s1_readdata;
  internal_clock_crossing_0_m1_requests_gpio1_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(7 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("01000000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --gpio1_s1_arb_share_counter set values, which is an e_mux
  gpio1_s1_arb_share_set_values <= std_logic'('1');
  --gpio1_s1_non_bursting_master_requests mux, which is an e_mux
  gpio1_s1_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_gpio1_s1;
  --gpio1_s1_any_bursting_master_saved_grant mux, which is an e_mux
  gpio1_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --gpio1_s1_arb_share_counter_next_value assignment, which is an e_assign
  gpio1_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gpio1_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpio1_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gpio1_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpio1_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gpio1_s1_allgrants all slave grants, which is an e_mux
  gpio1_s1_allgrants <= gpio1_s1_grant_vector;
  --gpio1_s1_end_xfer assignment, which is an e_assign
  gpio1_s1_end_xfer <= NOT ((gpio1_s1_waits_for_read OR gpio1_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_gpio1_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gpio1_s1 <= gpio1_s1_end_xfer AND (((NOT gpio1_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gpio1_s1_arb_share_counter arbitration counter enable, which is an e_assign
  gpio1_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gpio1_s1 AND gpio1_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_gpio1_s1 AND NOT gpio1_s1_non_bursting_master_requests));
  --gpio1_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpio1_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gpio1_s1_arb_counter_enable) = '1' then 
        gpio1_s1_arb_share_counter <= gpio1_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpio1_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpio1_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gpio1_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_gpio1_s1)) OR ((end_xfer_arb_share_counter_term_gpio1_s1 AND NOT gpio1_s1_non_bursting_master_requests)))) = '1' then 
        gpio1_s1_slavearbiterlockenable <= gpio1_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 gpio1/s1 arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= gpio1_s1_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --gpio1_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gpio1_s1_slavearbiterlockenable2 <= gpio1_s1_arb_share_counter_next_value;
  --clock_crossing_0/m1 gpio1/s1 arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= gpio1_s1_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --gpio1_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  gpio1_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_gpio1_s1 <= internal_clock_crossing_0_m1_requests_gpio1_s1 AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_gpio1_s1, which is an e_mux
  clock_crossing_0_m1_read_data_valid_gpio1_s1 <= (internal_clock_crossing_0_m1_granted_gpio1_s1 AND clock_crossing_0_m1_read) AND NOT gpio1_s1_waits_for_read;
  --gpio1_s1_writedata mux, which is an e_mux
  gpio1_s1_writedata <= clock_crossing_0_m1_writedata (7 DOWNTO 0);
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_gpio1_s1 <= internal_clock_crossing_0_m1_qualified_request_gpio1_s1;
  --clock_crossing_0/m1 saved-grant gpio1/s1, which is an e_assign
  clock_crossing_0_m1_saved_grant_gpio1_s1 <= internal_clock_crossing_0_m1_requests_gpio1_s1;
  --allow new arb cycle for gpio1/s1, which is an e_assign
  gpio1_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gpio1_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gpio1_s1_master_qreq_vector <= std_logic'('1');
  --gpio1_s1_reset_n assignment, which is an e_assign
  gpio1_s1_reset_n <= reset_n;
  gpio1_s1_chipselect <= internal_clock_crossing_0_m1_granted_gpio1_s1;
  --gpio1_s1_firsttransfer first transaction, which is an e_assign
  gpio1_s1_firsttransfer <= A_WE_StdLogic((std_logic'(gpio1_s1_begins_xfer) = '1'), gpio1_s1_unreg_firsttransfer, gpio1_s1_reg_firsttransfer);
  --gpio1_s1_unreg_firsttransfer first transaction, which is an e_assign
  gpio1_s1_unreg_firsttransfer <= NOT ((gpio1_s1_slavearbiterlockenable AND gpio1_s1_any_continuerequest));
  --gpio1_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpio1_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gpio1_s1_begins_xfer) = '1' then 
        gpio1_s1_reg_firsttransfer <= gpio1_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gpio1_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gpio1_s1_beginbursttransfer_internal <= gpio1_s1_begins_xfer;
  --~gpio1_s1_write_n assignment, which is an e_mux
  gpio1_s1_write_n <= NOT ((((internal_clock_crossing_0_m1_granted_gpio1_s1 AND clock_crossing_0_m1_write)) AND gpio1_s1_pretend_byte_enable));
  --gpio1_s1_address mux, which is an e_mux
  gpio1_s1_address <= clock_crossing_0_m1_nativeaddress (2 DOWNTO 0);
  --d1_gpio1_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gpio1_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gpio1_s1_end_xfer <= gpio1_s1_end_xfer;
    end if;

  end process;

  --gpio1_s1_waits_for_read in a cycle, which is an e_mux
  gpio1_s1_waits_for_read <= gpio1_s1_in_a_read_cycle AND gpio1_s1_begins_xfer;
  --gpio1_s1_in_a_read_cycle assignment, which is an e_assign
  gpio1_s1_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_gpio1_s1 AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gpio1_s1_in_a_read_cycle;
  --gpio1_s1_waits_for_write in a cycle, which is an e_mux
  gpio1_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpio1_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --gpio1_s1_in_a_write_cycle assignment, which is an e_assign
  gpio1_s1_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_gpio1_s1 AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gpio1_s1_in_a_write_cycle;
  wait_for_gpio1_s1_counter <= std_logic'('0');
  --gpio1_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  gpio1_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_clock_crossing_0_m1_granted_gpio1_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (clock_crossing_0_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_gpio1_s1 <= internal_clock_crossing_0_m1_granted_gpio1_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_gpio1_s1 <= internal_clock_crossing_0_m1_qualified_request_gpio1_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_gpio1_s1 <= internal_clock_crossing_0_m1_requests_gpio1_s1;
--synthesis translate_off
    --gpio1/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpio2_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal gpio2_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_m1_granted_gpio2_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_gpio2_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_gpio2_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_gpio2_s1 : OUT STD_LOGIC;
                 signal d1_gpio2_s1_end_xfer : OUT STD_LOGIC;
                 signal gpio2_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal gpio2_s1_chipselect : OUT STD_LOGIC;
                 signal gpio2_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gpio2_s1_reset_n : OUT STD_LOGIC;
                 signal gpio2_s1_write_n : OUT STD_LOGIC;
                 signal gpio2_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity gpio2_s1_arbitrator;


architecture europa of gpio2_s1_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_gpio2_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_gpio2_s1 :  STD_LOGIC;
                signal gpio2_s1_allgrants :  STD_LOGIC;
                signal gpio2_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal gpio2_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal gpio2_s1_any_continuerequest :  STD_LOGIC;
                signal gpio2_s1_arb_counter_enable :  STD_LOGIC;
                signal gpio2_s1_arb_share_counter :  STD_LOGIC;
                signal gpio2_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal gpio2_s1_arb_share_set_values :  STD_LOGIC;
                signal gpio2_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal gpio2_s1_begins_xfer :  STD_LOGIC;
                signal gpio2_s1_end_xfer :  STD_LOGIC;
                signal gpio2_s1_firsttransfer :  STD_LOGIC;
                signal gpio2_s1_grant_vector :  STD_LOGIC;
                signal gpio2_s1_in_a_read_cycle :  STD_LOGIC;
                signal gpio2_s1_in_a_write_cycle :  STD_LOGIC;
                signal gpio2_s1_master_qreq_vector :  STD_LOGIC;
                signal gpio2_s1_non_bursting_master_requests :  STD_LOGIC;
                signal gpio2_s1_pretend_byte_enable :  STD_LOGIC;
                signal gpio2_s1_reg_firsttransfer :  STD_LOGIC;
                signal gpio2_s1_slavearbiterlockenable :  STD_LOGIC;
                signal gpio2_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal gpio2_s1_unreg_firsttransfer :  STD_LOGIC;
                signal gpio2_s1_waits_for_read :  STD_LOGIC;
                signal gpio2_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_gpio2_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_gpio2_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_gpio2_s1 :  STD_LOGIC;
                signal wait_for_gpio2_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT gpio2_s1_end_xfer;
    end if;

  end process;

  gpio2_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_gpio2_s1);
  --assign gpio2_s1_readdata_from_sa = gpio2_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  gpio2_s1_readdata_from_sa <= gpio2_s1_readdata;
  internal_clock_crossing_0_m1_requests_gpio2_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(7 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("11000000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --gpio2_s1_arb_share_counter set values, which is an e_mux
  gpio2_s1_arb_share_set_values <= std_logic'('1');
  --gpio2_s1_non_bursting_master_requests mux, which is an e_mux
  gpio2_s1_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_gpio2_s1;
  --gpio2_s1_any_bursting_master_saved_grant mux, which is an e_mux
  gpio2_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --gpio2_s1_arb_share_counter_next_value assignment, which is an e_assign
  gpio2_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(gpio2_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpio2_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(gpio2_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpio2_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --gpio2_s1_allgrants all slave grants, which is an e_mux
  gpio2_s1_allgrants <= gpio2_s1_grant_vector;
  --gpio2_s1_end_xfer assignment, which is an e_assign
  gpio2_s1_end_xfer <= NOT ((gpio2_s1_waits_for_read OR gpio2_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_gpio2_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_gpio2_s1 <= gpio2_s1_end_xfer AND (((NOT gpio2_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --gpio2_s1_arb_share_counter arbitration counter enable, which is an e_assign
  gpio2_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_gpio2_s1 AND gpio2_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_gpio2_s1 AND NOT gpio2_s1_non_bursting_master_requests));
  --gpio2_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpio2_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(gpio2_s1_arb_counter_enable) = '1' then 
        gpio2_s1_arb_share_counter <= gpio2_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpio2_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpio2_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((gpio2_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_gpio2_s1)) OR ((end_xfer_arb_share_counter_term_gpio2_s1 AND NOT gpio2_s1_non_bursting_master_requests)))) = '1' then 
        gpio2_s1_slavearbiterlockenable <= gpio2_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 gpio2/s1 arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= gpio2_s1_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --gpio2_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  gpio2_s1_slavearbiterlockenable2 <= gpio2_s1_arb_share_counter_next_value;
  --clock_crossing_0/m1 gpio2/s1 arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= gpio2_s1_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --gpio2_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  gpio2_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_gpio2_s1 <= internal_clock_crossing_0_m1_requests_gpio2_s1 AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_gpio2_s1, which is an e_mux
  clock_crossing_0_m1_read_data_valid_gpio2_s1 <= (internal_clock_crossing_0_m1_granted_gpio2_s1 AND clock_crossing_0_m1_read) AND NOT gpio2_s1_waits_for_read;
  --gpio2_s1_writedata mux, which is an e_mux
  gpio2_s1_writedata <= clock_crossing_0_m1_writedata (7 DOWNTO 0);
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_gpio2_s1 <= internal_clock_crossing_0_m1_qualified_request_gpio2_s1;
  --clock_crossing_0/m1 saved-grant gpio2/s1, which is an e_assign
  clock_crossing_0_m1_saved_grant_gpio2_s1 <= internal_clock_crossing_0_m1_requests_gpio2_s1;
  --allow new arb cycle for gpio2/s1, which is an e_assign
  gpio2_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  gpio2_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  gpio2_s1_master_qreq_vector <= std_logic'('1');
  --gpio2_s1_reset_n assignment, which is an e_assign
  gpio2_s1_reset_n <= reset_n;
  gpio2_s1_chipselect <= internal_clock_crossing_0_m1_granted_gpio2_s1;
  --gpio2_s1_firsttransfer first transaction, which is an e_assign
  gpio2_s1_firsttransfer <= A_WE_StdLogic((std_logic'(gpio2_s1_begins_xfer) = '1'), gpio2_s1_unreg_firsttransfer, gpio2_s1_reg_firsttransfer);
  --gpio2_s1_unreg_firsttransfer first transaction, which is an e_assign
  gpio2_s1_unreg_firsttransfer <= NOT ((gpio2_s1_slavearbiterlockenable AND gpio2_s1_any_continuerequest));
  --gpio2_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpio2_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(gpio2_s1_begins_xfer) = '1' then 
        gpio2_s1_reg_firsttransfer <= gpio2_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --gpio2_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  gpio2_s1_beginbursttransfer_internal <= gpio2_s1_begins_xfer;
  --~gpio2_s1_write_n assignment, which is an e_mux
  gpio2_s1_write_n <= NOT ((((internal_clock_crossing_0_m1_granted_gpio2_s1 AND clock_crossing_0_m1_write)) AND gpio2_s1_pretend_byte_enable));
  --gpio2_s1_address mux, which is an e_mux
  gpio2_s1_address <= clock_crossing_0_m1_nativeaddress (1 DOWNTO 0);
  --d1_gpio2_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_gpio2_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_gpio2_s1_end_xfer <= gpio2_s1_end_xfer;
    end if;

  end process;

  --gpio2_s1_waits_for_read in a cycle, which is an e_mux
  gpio2_s1_waits_for_read <= gpio2_s1_in_a_read_cycle AND gpio2_s1_begins_xfer;
  --gpio2_s1_in_a_read_cycle assignment, which is an e_assign
  gpio2_s1_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_gpio2_s1 AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= gpio2_s1_in_a_read_cycle;
  --gpio2_s1_waits_for_write in a cycle, which is an e_mux
  gpio2_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(gpio2_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --gpio2_s1_in_a_write_cycle assignment, which is an e_assign
  gpio2_s1_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_gpio2_s1 AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= gpio2_s1_in_a_write_cycle;
  wait_for_gpio2_s1_counter <= std_logic'('0');
  --gpio2_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  gpio2_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_clock_crossing_0_m1_granted_gpio2_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (clock_crossing_0_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_gpio2_s1 <= internal_clock_crossing_0_m1_granted_gpio2_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_gpio2_s1 <= internal_clock_crossing_0_m1_qualified_request_gpio2_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_gpio2_s1 <= internal_clock_crossing_0_m1_requests_gpio2_s1;
--synthesis translate_off
    --gpio2/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity high_res_timer_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal high_res_timer_s1_irq : IN STD_LOGIC;
                 signal high_res_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_m1_granted_high_res_timer_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_high_res_timer_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_high_res_timer_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_high_res_timer_s1 : OUT STD_LOGIC;
                 signal d1_high_res_timer_s1_end_xfer : OUT STD_LOGIC;
                 signal high_res_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal high_res_timer_s1_chipselect : OUT STD_LOGIC;
                 signal high_res_timer_s1_irq_from_sa : OUT STD_LOGIC;
                 signal high_res_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal high_res_timer_s1_reset_n : OUT STD_LOGIC;
                 signal high_res_timer_s1_write_n : OUT STD_LOGIC;
                 signal high_res_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity high_res_timer_s1_arbitrator;


architecture europa of high_res_timer_s1_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_high_res_timer_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_high_res_timer_s1 :  STD_LOGIC;
                signal high_res_timer_s1_allgrants :  STD_LOGIC;
                signal high_res_timer_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal high_res_timer_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal high_res_timer_s1_any_continuerequest :  STD_LOGIC;
                signal high_res_timer_s1_arb_counter_enable :  STD_LOGIC;
                signal high_res_timer_s1_arb_share_counter :  STD_LOGIC;
                signal high_res_timer_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal high_res_timer_s1_arb_share_set_values :  STD_LOGIC;
                signal high_res_timer_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal high_res_timer_s1_begins_xfer :  STD_LOGIC;
                signal high_res_timer_s1_end_xfer :  STD_LOGIC;
                signal high_res_timer_s1_firsttransfer :  STD_LOGIC;
                signal high_res_timer_s1_grant_vector :  STD_LOGIC;
                signal high_res_timer_s1_in_a_read_cycle :  STD_LOGIC;
                signal high_res_timer_s1_in_a_write_cycle :  STD_LOGIC;
                signal high_res_timer_s1_master_qreq_vector :  STD_LOGIC;
                signal high_res_timer_s1_non_bursting_master_requests :  STD_LOGIC;
                signal high_res_timer_s1_reg_firsttransfer :  STD_LOGIC;
                signal high_res_timer_s1_slavearbiterlockenable :  STD_LOGIC;
                signal high_res_timer_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal high_res_timer_s1_unreg_firsttransfer :  STD_LOGIC;
                signal high_res_timer_s1_waits_for_read :  STD_LOGIC;
                signal high_res_timer_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_high_res_timer_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_high_res_timer_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_high_res_timer_s1 :  STD_LOGIC;
                signal wait_for_high_res_timer_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT high_res_timer_s1_end_xfer;
    end if;

  end process;

  high_res_timer_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_high_res_timer_s1);
  --assign high_res_timer_s1_readdata_from_sa = high_res_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  high_res_timer_s1_readdata_from_sa <= high_res_timer_s1_readdata;
  internal_clock_crossing_0_m1_requests_high_res_timer_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(7 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("00100000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --high_res_timer_s1_arb_share_counter set values, which is an e_mux
  high_res_timer_s1_arb_share_set_values <= std_logic'('1');
  --high_res_timer_s1_non_bursting_master_requests mux, which is an e_mux
  high_res_timer_s1_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_high_res_timer_s1;
  --high_res_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  high_res_timer_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --high_res_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  high_res_timer_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(high_res_timer_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(high_res_timer_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(high_res_timer_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(high_res_timer_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --high_res_timer_s1_allgrants all slave grants, which is an e_mux
  high_res_timer_s1_allgrants <= high_res_timer_s1_grant_vector;
  --high_res_timer_s1_end_xfer assignment, which is an e_assign
  high_res_timer_s1_end_xfer <= NOT ((high_res_timer_s1_waits_for_read OR high_res_timer_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_high_res_timer_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_high_res_timer_s1 <= high_res_timer_s1_end_xfer AND (((NOT high_res_timer_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --high_res_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  high_res_timer_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_high_res_timer_s1 AND high_res_timer_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_high_res_timer_s1 AND NOT high_res_timer_s1_non_bursting_master_requests));
  --high_res_timer_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      high_res_timer_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(high_res_timer_s1_arb_counter_enable) = '1' then 
        high_res_timer_s1_arb_share_counter <= high_res_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --high_res_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      high_res_timer_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((high_res_timer_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_high_res_timer_s1)) OR ((end_xfer_arb_share_counter_term_high_res_timer_s1 AND NOT high_res_timer_s1_non_bursting_master_requests)))) = '1' then 
        high_res_timer_s1_slavearbiterlockenable <= high_res_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 high_res_timer/s1 arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= high_res_timer_s1_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --high_res_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  high_res_timer_s1_slavearbiterlockenable2 <= high_res_timer_s1_arb_share_counter_next_value;
  --clock_crossing_0/m1 high_res_timer/s1 arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= high_res_timer_s1_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --high_res_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  high_res_timer_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_high_res_timer_s1 <= internal_clock_crossing_0_m1_requests_high_res_timer_s1 AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_high_res_timer_s1, which is an e_mux
  clock_crossing_0_m1_read_data_valid_high_res_timer_s1 <= (internal_clock_crossing_0_m1_granted_high_res_timer_s1 AND clock_crossing_0_m1_read) AND NOT high_res_timer_s1_waits_for_read;
  --high_res_timer_s1_writedata mux, which is an e_mux
  high_res_timer_s1_writedata <= clock_crossing_0_m1_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_high_res_timer_s1 <= internal_clock_crossing_0_m1_qualified_request_high_res_timer_s1;
  --clock_crossing_0/m1 saved-grant high_res_timer/s1, which is an e_assign
  clock_crossing_0_m1_saved_grant_high_res_timer_s1 <= internal_clock_crossing_0_m1_requests_high_res_timer_s1;
  --allow new arb cycle for high_res_timer/s1, which is an e_assign
  high_res_timer_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  high_res_timer_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  high_res_timer_s1_master_qreq_vector <= std_logic'('1');
  --high_res_timer_s1_reset_n assignment, which is an e_assign
  high_res_timer_s1_reset_n <= reset_n;
  high_res_timer_s1_chipselect <= internal_clock_crossing_0_m1_granted_high_res_timer_s1;
  --high_res_timer_s1_firsttransfer first transaction, which is an e_assign
  high_res_timer_s1_firsttransfer <= A_WE_StdLogic((std_logic'(high_res_timer_s1_begins_xfer) = '1'), high_res_timer_s1_unreg_firsttransfer, high_res_timer_s1_reg_firsttransfer);
  --high_res_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  high_res_timer_s1_unreg_firsttransfer <= NOT ((high_res_timer_s1_slavearbiterlockenable AND high_res_timer_s1_any_continuerequest));
  --high_res_timer_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      high_res_timer_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(high_res_timer_s1_begins_xfer) = '1' then 
        high_res_timer_s1_reg_firsttransfer <= high_res_timer_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --high_res_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  high_res_timer_s1_beginbursttransfer_internal <= high_res_timer_s1_begins_xfer;
  --~high_res_timer_s1_write_n assignment, which is an e_mux
  high_res_timer_s1_write_n <= NOT ((internal_clock_crossing_0_m1_granted_high_res_timer_s1 AND clock_crossing_0_m1_write));
  --high_res_timer_s1_address mux, which is an e_mux
  high_res_timer_s1_address <= clock_crossing_0_m1_nativeaddress (2 DOWNTO 0);
  --d1_high_res_timer_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_high_res_timer_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_high_res_timer_s1_end_xfer <= high_res_timer_s1_end_xfer;
    end if;

  end process;

  --high_res_timer_s1_waits_for_read in a cycle, which is an e_mux
  high_res_timer_s1_waits_for_read <= high_res_timer_s1_in_a_read_cycle AND high_res_timer_s1_begins_xfer;
  --high_res_timer_s1_in_a_read_cycle assignment, which is an e_assign
  high_res_timer_s1_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_high_res_timer_s1 AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= high_res_timer_s1_in_a_read_cycle;
  --high_res_timer_s1_waits_for_write in a cycle, which is an e_mux
  high_res_timer_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(high_res_timer_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --high_res_timer_s1_in_a_write_cycle assignment, which is an e_assign
  high_res_timer_s1_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_high_res_timer_s1 AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= high_res_timer_s1_in_a_write_cycle;
  wait_for_high_res_timer_s1_counter <= std_logic'('0');
  --assign high_res_timer_s1_irq_from_sa = high_res_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  high_res_timer_s1_irq_from_sa <= high_res_timer_s1_irq;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_high_res_timer_s1 <= internal_clock_crossing_0_m1_granted_high_res_timer_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_high_res_timer_s1 <= internal_clock_crossing_0_m1_qualified_request_high_res_timer_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_high_res_timer_s1 <= internal_clock_crossing_0_m1_requests_high_res_timer_s1;
--synthesis translate_off
    --high_res_timer/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity jtag_uart_avalon_jtag_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity jtag_uart_avalon_jtag_slave_arbitrator;


architecture europa of jtag_uart_avalon_jtag_slave_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allgrants :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_continuerequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_counter_enable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_counter :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_set_values :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_begins_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_grant_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_read_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_write_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_master_qreq_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_non_bursting_master_requests :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_unreg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_read :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_write :  STD_LOGIC;
                signal wait_for_jtag_uart_avalon_jtag_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  jtag_uart_avalon_jtag_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave);
  --assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readdata_from_sa <= jtag_uart_avalon_jtag_slave_readdata;
  internal_clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(7 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("11010000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_dataavailable_from_sa <= jtag_uart_avalon_jtag_slave_dataavailable;
  --assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readyfordata_from_sa <= jtag_uart_avalon_jtag_slave_readyfordata;
  --assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= jtag_uart_avalon_jtag_slave_waitrequest;
  --jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  jtag_uart_avalon_jtag_slave_arb_share_set_values <= std_logic'('1');
  --jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(jtag_uart_avalon_jtag_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_avalon_jtag_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(jtag_uart_avalon_jtag_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_avalon_jtag_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  jtag_uart_avalon_jtag_slave_allgrants <= jtag_uart_avalon_jtag_slave_grant_vector;
  --jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_end_xfer <= NOT ((jtag_uart_avalon_jtag_slave_waits_for_read OR jtag_uart_avalon_jtag_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave <= jtag_uart_avalon_jtag_slave_end_xfer AND (((NOT jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND jtag_uart_avalon_jtag_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests));
  --jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_arb_counter_enable) = '1' then 
        jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((jtag_uart_avalon_jtag_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests)))) = '1' then 
        jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
  --clock_crossing_0/m1 jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  jtag_uart_avalon_jtag_slave_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave <= internal_clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave, which is an e_mux
  clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave <= (internal_clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave AND clock_crossing_0_m1_read) AND NOT jtag_uart_avalon_jtag_slave_waits_for_read;
  --jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_writedata <= clock_crossing_0_m1_writedata;
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave <= internal_clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  --clock_crossing_0/m1 saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  clock_crossing_0_m1_saved_grant_jtag_uart_avalon_jtag_slave <= internal_clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave;
  --allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  jtag_uart_avalon_jtag_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  jtag_uart_avalon_jtag_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  jtag_uart_avalon_jtag_slave_master_qreq_vector <= std_logic'('1');
  --jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_reset_n <= reset_n;
  jtag_uart_avalon_jtag_slave_chipselect <= internal_clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_firsttransfer <= A_WE_StdLogic((std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1'), jtag_uart_avalon_jtag_slave_unreg_firsttransfer, jtag_uart_avalon_jtag_slave_reg_firsttransfer);
  --jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_unreg_firsttransfer <= NOT ((jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND jtag_uart_avalon_jtag_slave_any_continuerequest));
  --jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1' then 
        jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  jtag_uart_avalon_jtag_slave_beginbursttransfer_internal <= jtag_uart_avalon_jtag_slave_begins_xfer;
  --~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_read_n <= NOT ((internal_clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave AND clock_crossing_0_m1_read));
  --~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_write_n <= NOT ((internal_clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave AND clock_crossing_0_m1_write));
  --jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_address <= clock_crossing_0_m1_nativeaddress(0);
  --d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_read <= jtag_uart_avalon_jtag_slave_in_a_read_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  --jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_write <= jtag_uart_avalon_jtag_slave_in_a_write_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wait_for_jtag_uart_avalon_jtag_slave_counter <= std_logic'('0');
  --assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_irq_from_sa <= jtag_uart_avalon_jtag_slave_irq;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave <= internal_clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave <= internal_clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave <= internal_clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
--synthesis translate_off
    --jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity led_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal led_pio_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_m1_granted_led_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_led_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_led_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_led_pio_s1 : OUT STD_LOGIC;
                 signal d1_led_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal led_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal led_pio_s1_chipselect : OUT STD_LOGIC;
                 signal led_pio_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal led_pio_s1_reset_n : OUT STD_LOGIC;
                 signal led_pio_s1_write_n : OUT STD_LOGIC;
                 signal led_pio_s1_writedata : OUT STD_LOGIC
              );
end entity led_pio_s1_arbitrator;


architecture europa of led_pio_s1_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_led_pio_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_led_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_led_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_led_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_led_pio_s1 :  STD_LOGIC;
                signal led_pio_s1_allgrants :  STD_LOGIC;
                signal led_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal led_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal led_pio_s1_any_continuerequest :  STD_LOGIC;
                signal led_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal led_pio_s1_arb_share_counter :  STD_LOGIC;
                signal led_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal led_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal led_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal led_pio_s1_begins_xfer :  STD_LOGIC;
                signal led_pio_s1_end_xfer :  STD_LOGIC;
                signal led_pio_s1_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_grant_vector :  STD_LOGIC;
                signal led_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal led_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal led_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal led_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal led_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal led_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal led_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_waits_for_read :  STD_LOGIC;
                signal led_pio_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_led_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT led_pio_s1_end_xfer;
    end if;

  end process;

  led_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_led_pio_s1);
  --assign led_pio_s1_readdata_from_sa = led_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  led_pio_s1_readdata_from_sa <= led_pio_s1_readdata;
  internal_clock_crossing_0_m1_requests_led_pio_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(7 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10100000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --led_pio_s1_arb_share_counter set values, which is an e_mux
  led_pio_s1_arb_share_set_values <= std_logic'('1');
  --led_pio_s1_non_bursting_master_requests mux, which is an e_mux
  led_pio_s1_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_led_pio_s1;
  --led_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  led_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --led_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  led_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(led_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(led_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --led_pio_s1_allgrants all slave grants, which is an e_mux
  led_pio_s1_allgrants <= led_pio_s1_grant_vector;
  --led_pio_s1_end_xfer assignment, which is an e_assign
  led_pio_s1_end_xfer <= NOT ((led_pio_s1_waits_for_read OR led_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_led_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_led_pio_s1 <= led_pio_s1_end_xfer AND (((NOT led_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --led_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  led_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_led_pio_s1 AND led_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_led_pio_s1 AND NOT led_pio_s1_non_bursting_master_requests));
  --led_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(led_pio_s1_arb_counter_enable) = '1' then 
        led_pio_s1_arb_share_counter <= led_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --led_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((led_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_led_pio_s1)) OR ((end_xfer_arb_share_counter_term_led_pio_s1 AND NOT led_pio_s1_non_bursting_master_requests)))) = '1' then 
        led_pio_s1_slavearbiterlockenable <= led_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 led_pio/s1 arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= led_pio_s1_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --led_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  led_pio_s1_slavearbiterlockenable2 <= led_pio_s1_arb_share_counter_next_value;
  --clock_crossing_0/m1 led_pio/s1 arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= led_pio_s1_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --led_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  led_pio_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_led_pio_s1 <= internal_clock_crossing_0_m1_requests_led_pio_s1 AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_led_pio_s1, which is an e_mux
  clock_crossing_0_m1_read_data_valid_led_pio_s1 <= (internal_clock_crossing_0_m1_granted_led_pio_s1 AND clock_crossing_0_m1_read) AND NOT led_pio_s1_waits_for_read;
  --led_pio_s1_writedata mux, which is an e_mux
  led_pio_s1_writedata <= clock_crossing_0_m1_writedata(0);
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_led_pio_s1 <= internal_clock_crossing_0_m1_qualified_request_led_pio_s1;
  --clock_crossing_0/m1 saved-grant led_pio/s1, which is an e_assign
  clock_crossing_0_m1_saved_grant_led_pio_s1 <= internal_clock_crossing_0_m1_requests_led_pio_s1;
  --allow new arb cycle for led_pio/s1, which is an e_assign
  led_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  led_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  led_pio_s1_master_qreq_vector <= std_logic'('1');
  --led_pio_s1_reset_n assignment, which is an e_assign
  led_pio_s1_reset_n <= reset_n;
  led_pio_s1_chipselect <= internal_clock_crossing_0_m1_granted_led_pio_s1;
  --led_pio_s1_firsttransfer first transaction, which is an e_assign
  led_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(led_pio_s1_begins_xfer) = '1'), led_pio_s1_unreg_firsttransfer, led_pio_s1_reg_firsttransfer);
  --led_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  led_pio_s1_unreg_firsttransfer <= NOT ((led_pio_s1_slavearbiterlockenable AND led_pio_s1_any_continuerequest));
  --led_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(led_pio_s1_begins_xfer) = '1' then 
        led_pio_s1_reg_firsttransfer <= led_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --led_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  led_pio_s1_beginbursttransfer_internal <= led_pio_s1_begins_xfer;
  --~led_pio_s1_write_n assignment, which is an e_mux
  led_pio_s1_write_n <= NOT ((internal_clock_crossing_0_m1_granted_led_pio_s1 AND clock_crossing_0_m1_write));
  --led_pio_s1_address mux, which is an e_mux
  led_pio_s1_address <= clock_crossing_0_m1_nativeaddress (1 DOWNTO 0);
  --d1_led_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_led_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_led_pio_s1_end_xfer <= led_pio_s1_end_xfer;
    end if;

  end process;

  --led_pio_s1_waits_for_read in a cycle, which is an e_mux
  led_pio_s1_waits_for_read <= led_pio_s1_in_a_read_cycle AND led_pio_s1_begins_xfer;
  --led_pio_s1_in_a_read_cycle assignment, which is an e_assign
  led_pio_s1_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_led_pio_s1 AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= led_pio_s1_in_a_read_cycle;
  --led_pio_s1_waits_for_write in a cycle, which is an e_mux
  led_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --led_pio_s1_in_a_write_cycle assignment, which is an e_assign
  led_pio_s1_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_led_pio_s1 AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= led_pio_s1_in_a_write_cycle;
  wait_for_led_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_led_pio_s1 <= internal_clock_crossing_0_m1_granted_led_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_led_pio_s1 <= internal_clock_crossing_0_m1_qualified_request_led_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_led_pio_s1 <= internal_clock_crossing_0_m1_requests_led_pio_s1;
--synthesis translate_off
    --led_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity onchip_memory_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_0_data_master_read : IN STD_LOGIC;
                 signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                 signal cpu_0_data_master_write : IN STD_LOGIC;
                 signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_0_instruction_master_read : IN STD_LOGIC;
                 signal onchip_memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_0_data_master_granted_onchip_memory_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_qualified_request_onchip_memory_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_read_data_valid_onchip_memory_s1 : OUT STD_LOGIC;
                 signal cpu_0_data_master_requests_onchip_memory_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_granted_onchip_memory_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_qualified_request_onchip_memory_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_read_data_valid_onchip_memory_s1 : OUT STD_LOGIC;
                 signal cpu_0_instruction_master_requests_onchip_memory_s1 : OUT STD_LOGIC;
                 signal d1_onchip_memory_s1_end_xfer : OUT STD_LOGIC;
                 signal onchip_memory_s1_address : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal onchip_memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal onchip_memory_s1_chipselect : OUT STD_LOGIC;
                 signal onchip_memory_s1_clken : OUT STD_LOGIC;
                 signal onchip_memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal onchip_memory_s1_reset : OUT STD_LOGIC;
                 signal onchip_memory_s1_write : OUT STD_LOGIC;
                 signal onchip_memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal registered_cpu_0_data_master_read_data_valid_onchip_memory_s1 : OUT STD_LOGIC
              );
end entity onchip_memory_s1_arbitrator;


architecture europa of onchip_memory_s1_arbitrator is
                signal cpu_0_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_data_master_continuerequest :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register_in :  STD_LOGIC;
                signal cpu_0_data_master_saved_grant_onchip_memory_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_0_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_0_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register_in :  STD_LOGIC;
                signal cpu_0_instruction_master_saved_grant_onchip_memory_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_onchip_memory_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_0_data_master_granted_onchip_memory_s1 :  STD_LOGIC;
                signal internal_cpu_0_data_master_qualified_request_onchip_memory_s1 :  STD_LOGIC;
                signal internal_cpu_0_data_master_requests_onchip_memory_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_granted_onchip_memory_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_qualified_request_onchip_memory_s1 :  STD_LOGIC;
                signal internal_cpu_0_instruction_master_requests_onchip_memory_s1 :  STD_LOGIC;
                signal last_cycle_cpu_0_data_master_granted_slave_onchip_memory_s1 :  STD_LOGIC;
                signal last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory_s1 :  STD_LOGIC;
                signal onchip_memory_s1_allgrants :  STD_LOGIC;
                signal onchip_memory_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal onchip_memory_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal onchip_memory_s1_any_continuerequest :  STD_LOGIC;
                signal onchip_memory_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_s1_arb_counter_enable :  STD_LOGIC;
                signal onchip_memory_s1_arb_share_counter :  STD_LOGIC;
                signal onchip_memory_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal onchip_memory_s1_arb_share_set_values :  STD_LOGIC;
                signal onchip_memory_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal onchip_memory_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal onchip_memory_s1_begins_xfer :  STD_LOGIC;
                signal onchip_memory_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal onchip_memory_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_s1_end_xfer :  STD_LOGIC;
                signal onchip_memory_s1_firsttransfer :  STD_LOGIC;
                signal onchip_memory_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_s1_in_a_read_cycle :  STD_LOGIC;
                signal onchip_memory_s1_in_a_write_cycle :  STD_LOGIC;
                signal onchip_memory_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_s1_non_bursting_master_requests :  STD_LOGIC;
                signal onchip_memory_s1_reg_firsttransfer :  STD_LOGIC;
                signal onchip_memory_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_s1_slavearbiterlockenable :  STD_LOGIC;
                signal onchip_memory_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal onchip_memory_s1_unreg_firsttransfer :  STD_LOGIC;
                signal onchip_memory_s1_waits_for_read :  STD_LOGIC;
                signal onchip_memory_s1_waits_for_write :  STD_LOGIC;
                signal p1_cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register :  STD_LOGIC;
                signal p1_cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register :  STD_LOGIC;
                signal shifted_address_to_onchip_memory_s1_from_cpu_0_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal shifted_address_to_onchip_memory_s1_from_cpu_0_instruction_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_onchip_memory_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT onchip_memory_s1_end_xfer;
    end if;

  end process;

  onchip_memory_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpu_0_data_master_qualified_request_onchip_memory_s1 OR internal_cpu_0_instruction_master_qualified_request_onchip_memory_s1));
  --assign onchip_memory_s1_readdata_from_sa = onchip_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  onchip_memory_s1_readdata_from_sa <= onchip_memory_s1_readdata;
  internal_cpu_0_data_master_requests_onchip_memory_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_0_data_master_address_to_slave(27 DOWNTO 14) & std_logic_vector'("00000000000000")) = std_logic_vector'("1010000000000100000000000000")))) AND ((cpu_0_data_master_read OR cpu_0_data_master_write));
  --registered rdv signal_name registered_cpu_0_data_master_read_data_valid_onchip_memory_s1 assignment, which is an e_assign
  registered_cpu_0_data_master_read_data_valid_onchip_memory_s1 <= cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register_in;
  --onchip_memory_s1_arb_share_counter set values, which is an e_mux
  onchip_memory_s1_arb_share_set_values <= std_logic'('1');
  --onchip_memory_s1_non_bursting_master_requests mux, which is an e_mux
  onchip_memory_s1_non_bursting_master_requests <= ((internal_cpu_0_data_master_requests_onchip_memory_s1 OR internal_cpu_0_instruction_master_requests_onchip_memory_s1) OR internal_cpu_0_data_master_requests_onchip_memory_s1) OR internal_cpu_0_instruction_master_requests_onchip_memory_s1;
  --onchip_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  onchip_memory_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --onchip_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  onchip_memory_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(onchip_memory_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(onchip_memory_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(onchip_memory_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(onchip_memory_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --onchip_memory_s1_allgrants all slave grants, which is an e_mux
  onchip_memory_s1_allgrants <= (((or_reduce(onchip_memory_s1_grant_vector)) OR (or_reduce(onchip_memory_s1_grant_vector))) OR (or_reduce(onchip_memory_s1_grant_vector))) OR (or_reduce(onchip_memory_s1_grant_vector));
  --onchip_memory_s1_end_xfer assignment, which is an e_assign
  onchip_memory_s1_end_xfer <= NOT ((onchip_memory_s1_waits_for_read OR onchip_memory_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_onchip_memory_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_onchip_memory_s1 <= onchip_memory_s1_end_xfer AND (((NOT onchip_memory_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --onchip_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  onchip_memory_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_onchip_memory_s1 AND onchip_memory_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_onchip_memory_s1 AND NOT onchip_memory_s1_non_bursting_master_requests));
  --onchip_memory_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_memory_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(onchip_memory_s1_arb_counter_enable) = '1' then 
        onchip_memory_s1_arb_share_counter <= onchip_memory_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --onchip_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_memory_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(onchip_memory_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_onchip_memory_s1)) OR ((end_xfer_arb_share_counter_term_onchip_memory_s1 AND NOT onchip_memory_s1_non_bursting_master_requests)))) = '1' then 
        onchip_memory_s1_slavearbiterlockenable <= onchip_memory_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_0/data_master onchip_memory/s1 arbiterlock, which is an e_assign
  cpu_0_data_master_arbiterlock <= onchip_memory_s1_slavearbiterlockenable AND cpu_0_data_master_continuerequest;
  --onchip_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  onchip_memory_s1_slavearbiterlockenable2 <= onchip_memory_s1_arb_share_counter_next_value;
  --cpu_0/data_master onchip_memory/s1 arbiterlock2, which is an e_assign
  cpu_0_data_master_arbiterlock2 <= onchip_memory_s1_slavearbiterlockenable2 AND cpu_0_data_master_continuerequest;
  --cpu_0/instruction_master onchip_memory/s1 arbiterlock, which is an e_assign
  cpu_0_instruction_master_arbiterlock <= onchip_memory_s1_slavearbiterlockenable AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master onchip_memory/s1 arbiterlock2, which is an e_assign
  cpu_0_instruction_master_arbiterlock2 <= onchip_memory_s1_slavearbiterlockenable2 AND cpu_0_instruction_master_continuerequest;
  --cpu_0/instruction_master granted onchip_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_instruction_master_saved_grant_onchip_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((onchip_memory_s1_arbitration_holdoff_internal OR NOT internal_cpu_0_instruction_master_requests_onchip_memory_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory_s1))))));
    end if;

  end process;

  --cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  cpu_0_instruction_master_continuerequest <= last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory_s1 AND internal_cpu_0_instruction_master_requests_onchip_memory_s1;
  --onchip_memory_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  onchip_memory_s1_any_continuerequest <= cpu_0_instruction_master_continuerequest OR cpu_0_data_master_continuerequest;
  internal_cpu_0_data_master_qualified_request_onchip_memory_s1 <= internal_cpu_0_data_master_requests_onchip_memory_s1 AND NOT (((((cpu_0_data_master_read AND (cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register))) OR (((NOT cpu_0_data_master_waitrequest) AND cpu_0_data_master_write))) OR cpu_0_instruction_master_arbiterlock));
  --cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register_in <= ((internal_cpu_0_data_master_granted_onchip_memory_s1 AND cpu_0_data_master_read) AND NOT onchip_memory_s1_waits_for_read) AND NOT (cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register);
  --shift register p1 cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register) & A_ToStdLogicVector(cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register_in)));
  --cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register <= p1_cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_0_data_master_read_data_valid_onchip_memory_s1, which is an e_mux
  cpu_0_data_master_read_data_valid_onchip_memory_s1 <= cpu_0_data_master_read_data_valid_onchip_memory_s1_shift_register;
  --onchip_memory_s1_writedata mux, which is an e_mux
  onchip_memory_s1_writedata <= cpu_0_data_master_writedata;
  --mux onchip_memory_s1_clken, which is an e_mux
  onchip_memory_s1_clken <= std_logic'('1');
  internal_cpu_0_instruction_master_requests_onchip_memory_s1 <= ((to_std_logic(((Std_Logic_Vector'(cpu_0_instruction_master_address_to_slave(27 DOWNTO 14) & std_logic_vector'("00000000000000")) = std_logic_vector'("1010000000000100000000000000")))) AND (cpu_0_instruction_master_read))) AND cpu_0_instruction_master_read;
  --cpu_0/data_master granted onchip_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_0_data_master_granted_slave_onchip_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_0_data_master_granted_slave_onchip_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_0_data_master_saved_grant_onchip_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((onchip_memory_s1_arbitration_holdoff_internal OR NOT internal_cpu_0_data_master_requests_onchip_memory_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_0_data_master_granted_slave_onchip_memory_s1))))));
    end if;

  end process;

  --cpu_0_data_master_continuerequest continued request, which is an e_mux
  cpu_0_data_master_continuerequest <= last_cycle_cpu_0_data_master_granted_slave_onchip_memory_s1 AND internal_cpu_0_data_master_requests_onchip_memory_s1;
  internal_cpu_0_instruction_master_qualified_request_onchip_memory_s1 <= internal_cpu_0_instruction_master_requests_onchip_memory_s1 AND NOT ((((cpu_0_instruction_master_read AND (cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register))) OR cpu_0_data_master_arbiterlock));
  --cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register_in <= ((internal_cpu_0_instruction_master_granted_onchip_memory_s1 AND cpu_0_instruction_master_read) AND NOT onchip_memory_s1_waits_for_read) AND NOT (cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register);
  --shift register p1 cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register) & A_ToStdLogicVector(cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register_in)));
  --cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register <= p1_cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_0_instruction_master_read_data_valid_onchip_memory_s1, which is an e_mux
  cpu_0_instruction_master_read_data_valid_onchip_memory_s1 <= cpu_0_instruction_master_read_data_valid_onchip_memory_s1_shift_register;
  --allow new arb cycle for onchip_memory/s1, which is an e_assign
  onchip_memory_s1_allow_new_arb_cycle <= NOT cpu_0_data_master_arbiterlock AND NOT cpu_0_instruction_master_arbiterlock;
  --cpu_0/instruction_master assignment into master qualified-requests vector for onchip_memory/s1, which is an e_assign
  onchip_memory_s1_master_qreq_vector(0) <= internal_cpu_0_instruction_master_qualified_request_onchip_memory_s1;
  --cpu_0/instruction_master grant onchip_memory/s1, which is an e_assign
  internal_cpu_0_instruction_master_granted_onchip_memory_s1 <= onchip_memory_s1_grant_vector(0);
  --cpu_0/instruction_master saved-grant onchip_memory/s1, which is an e_assign
  cpu_0_instruction_master_saved_grant_onchip_memory_s1 <= onchip_memory_s1_arb_winner(0) AND internal_cpu_0_instruction_master_requests_onchip_memory_s1;
  --cpu_0/data_master assignment into master qualified-requests vector for onchip_memory/s1, which is an e_assign
  onchip_memory_s1_master_qreq_vector(1) <= internal_cpu_0_data_master_qualified_request_onchip_memory_s1;
  --cpu_0/data_master grant onchip_memory/s1, which is an e_assign
  internal_cpu_0_data_master_granted_onchip_memory_s1 <= onchip_memory_s1_grant_vector(1);
  --cpu_0/data_master saved-grant onchip_memory/s1, which is an e_assign
  cpu_0_data_master_saved_grant_onchip_memory_s1 <= onchip_memory_s1_arb_winner(1) AND internal_cpu_0_data_master_requests_onchip_memory_s1;
  --onchip_memory/s1 chosen-master double-vector, which is an e_assign
  onchip_memory_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((onchip_memory_s1_master_qreq_vector & onchip_memory_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT onchip_memory_s1_master_qreq_vector & NOT onchip_memory_s1_master_qreq_vector))) + (std_logic_vector'("000") & (onchip_memory_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  onchip_memory_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((onchip_memory_s1_allow_new_arb_cycle AND or_reduce(onchip_memory_s1_grant_vector)))) = '1'), onchip_memory_s1_grant_vector, onchip_memory_s1_saved_chosen_master_vector);
  --saved onchip_memory_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_memory_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(onchip_memory_s1_allow_new_arb_cycle) = '1' then 
        onchip_memory_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(onchip_memory_s1_grant_vector)) = '1'), onchip_memory_s1_grant_vector, onchip_memory_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  onchip_memory_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((onchip_memory_s1_chosen_master_double_vector(1) OR onchip_memory_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((onchip_memory_s1_chosen_master_double_vector(0) OR onchip_memory_s1_chosen_master_double_vector(2)))));
  --onchip_memory/s1 chosen master rotated left, which is an e_assign
  onchip_memory_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(onchip_memory_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(onchip_memory_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --onchip_memory/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_memory_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(onchip_memory_s1_grant_vector)) = '1' then 
        onchip_memory_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(onchip_memory_s1_end_xfer) = '1'), onchip_memory_s1_chosen_master_rot_left, onchip_memory_s1_grant_vector);
      end if;
    end if;

  end process;

  --~onchip_memory_s1_reset assignment, which is an e_assign
  onchip_memory_s1_reset <= NOT reset_n;
  onchip_memory_s1_chipselect <= internal_cpu_0_data_master_granted_onchip_memory_s1 OR internal_cpu_0_instruction_master_granted_onchip_memory_s1;
  --onchip_memory_s1_firsttransfer first transaction, which is an e_assign
  onchip_memory_s1_firsttransfer <= A_WE_StdLogic((std_logic'(onchip_memory_s1_begins_xfer) = '1'), onchip_memory_s1_unreg_firsttransfer, onchip_memory_s1_reg_firsttransfer);
  --onchip_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  onchip_memory_s1_unreg_firsttransfer <= NOT ((onchip_memory_s1_slavearbiterlockenable AND onchip_memory_s1_any_continuerequest));
  --onchip_memory_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_memory_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(onchip_memory_s1_begins_xfer) = '1' then 
        onchip_memory_s1_reg_firsttransfer <= onchip_memory_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --onchip_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  onchip_memory_s1_beginbursttransfer_internal <= onchip_memory_s1_begins_xfer;
  --onchip_memory_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  onchip_memory_s1_arbitration_holdoff_internal <= onchip_memory_s1_begins_xfer AND onchip_memory_s1_firsttransfer;
  --onchip_memory_s1_write assignment, which is an e_mux
  onchip_memory_s1_write <= internal_cpu_0_data_master_granted_onchip_memory_s1 AND cpu_0_data_master_write;
  shifted_address_to_onchip_memory_s1_from_cpu_0_data_master <= cpu_0_data_master_address_to_slave;
  --onchip_memory_s1_address mux, which is an e_mux
  onchip_memory_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_onchip_memory_s1)) = '1'), (A_SRL(shifted_address_to_onchip_memory_s1_from_cpu_0_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_onchip_memory_s1_from_cpu_0_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 12);
  shifted_address_to_onchip_memory_s1_from_cpu_0_instruction_master <= cpu_0_instruction_master_address_to_slave;
  --d1_onchip_memory_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_onchip_memory_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_onchip_memory_s1_end_xfer <= onchip_memory_s1_end_xfer;
    end if;

  end process;

  --onchip_memory_s1_waits_for_read in a cycle, which is an e_mux
  onchip_memory_s1_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(onchip_memory_s1_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --onchip_memory_s1_in_a_read_cycle assignment, which is an e_assign
  onchip_memory_s1_in_a_read_cycle <= ((internal_cpu_0_data_master_granted_onchip_memory_s1 AND cpu_0_data_master_read)) OR ((internal_cpu_0_instruction_master_granted_onchip_memory_s1 AND cpu_0_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= onchip_memory_s1_in_a_read_cycle;
  --onchip_memory_s1_waits_for_write in a cycle, which is an e_mux
  onchip_memory_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(onchip_memory_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --onchip_memory_s1_in_a_write_cycle assignment, which is an e_assign
  onchip_memory_s1_in_a_write_cycle <= internal_cpu_0_data_master_granted_onchip_memory_s1 AND cpu_0_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= onchip_memory_s1_in_a_write_cycle;
  wait_for_onchip_memory_s1_counter <= std_logic'('0');
  --onchip_memory_s1_byteenable byte enable port mux, which is an e_mux
  onchip_memory_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_0_data_master_granted_onchip_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_0_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_0_data_master_granted_onchip_memory_s1 <= internal_cpu_0_data_master_granted_onchip_memory_s1;
  --vhdl renameroo for output signals
  cpu_0_data_master_qualified_request_onchip_memory_s1 <= internal_cpu_0_data_master_qualified_request_onchip_memory_s1;
  --vhdl renameroo for output signals
  cpu_0_data_master_requests_onchip_memory_s1 <= internal_cpu_0_data_master_requests_onchip_memory_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_granted_onchip_memory_s1 <= internal_cpu_0_instruction_master_granted_onchip_memory_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_qualified_request_onchip_memory_s1 <= internal_cpu_0_instruction_master_qualified_request_onchip_memory_s1;
  --vhdl renameroo for output signals
  cpu_0_instruction_master_requests_onchip_memory_s1 <= internal_cpu_0_instruction_master_requests_onchip_memory_s1;
--synthesis translate_off
    --onchip_memory/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line50 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_data_master_granted_onchip_memory_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_0_instruction_master_granted_onchip_memory_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line50, now);
          write(write_line50, string'(": "));
          write(write_line50, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line50.all);
          deallocate (write_line50);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line51 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_data_master_saved_grant_onchip_memory_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_0_instruction_master_saved_grant_onchip_memory_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line51, now);
          write(write_line51, string'(": "));
          write(write_line51, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line51.all);
          deallocate (write_line51);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_flash_ssram_pipeline_bridge_m1_to_pipeline_bridge_before_tristate_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_flash_ssram_pipeline_bridge_m1_to_pipeline_bridge_before_tristate_s1_module;


architecture europa of rdv_fifo_for_flash_ssram_pipeline_bridge_m1_to_pipeline_bridge_before_tristate_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pipeline_bridge_before_tristate_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal flash_ssram_pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_debugaccess : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_s1_endofpacket : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_s1_readdatavalid : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pipeline_bridge_before_tristate_s1_end_xfer : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1 : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1_shift_register : OUT STD_LOGIC;
                 signal flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_s1_arbiterlock : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_arbiterlock2 : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_burstcount : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_s1_chipselect : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_debugaccess : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_s1_read : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_s1_reset_n : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_write : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity pipeline_bridge_before_tristate_s1_arbitrator;


architecture europa of pipeline_bridge_before_tristate_s1_arbitrator is
component rdv_fifo_for_flash_ssram_pipeline_bridge_m1_to_pipeline_bridge_before_tristate_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_flash_ssram_pipeline_bridge_m1_to_pipeline_bridge_before_tristate_s1_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_rdv_fifo_empty_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_rdv_fifo_output_from_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_saved_grant_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal internal_flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal internal_flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_before_tristate_s1_waitrequest_from_sa :  STD_LOGIC;
                signal module_input22 :  STD_LOGIC;
                signal module_input23 :  STD_LOGIC;
                signal module_input24 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_allgrants :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_any_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_arb_counter_enable :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_arb_share_counter :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_arb_share_set_values :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_begins_xfer :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_end_xfer :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_firsttransfer :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_grant_vector :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_in_a_read_cycle :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_in_a_write_cycle :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_master_qreq_vector :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_reg_firsttransfer :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_waits_for_read :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pipeline_bridge_before_tristate_s1_from_flash_ssram_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_pipeline_bridge_before_tristate_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pipeline_bridge_before_tristate_s1_end_xfer;
    end if;

  end process;

  pipeline_bridge_before_tristate_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1);
  --assign pipeline_bridge_before_tristate_s1_readdata_from_sa = pipeline_bridge_before_tristate_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pipeline_bridge_before_tristate_s1_readdata_from_sa <= pipeline_bridge_before_tristate_s1_readdata;
  internal_flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(flash_ssram_pipeline_bridge_m1_chipselect)))));
  --assign pipeline_bridge_before_tristate_s1_waitrequest_from_sa = pipeline_bridge_before_tristate_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_pipeline_bridge_before_tristate_s1_waitrequest_from_sa <= pipeline_bridge_before_tristate_s1_waitrequest;
  --assign pipeline_bridge_before_tristate_s1_readdatavalid_from_sa = pipeline_bridge_before_tristate_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  pipeline_bridge_before_tristate_s1_readdatavalid_from_sa <= pipeline_bridge_before_tristate_s1_readdatavalid;
  --pipeline_bridge_before_tristate_s1_arb_share_counter set values, which is an e_mux
  pipeline_bridge_before_tristate_s1_arb_share_set_values <= std_logic'('1');
  --pipeline_bridge_before_tristate_s1_non_bursting_master_requests mux, which is an e_mux
  pipeline_bridge_before_tristate_s1_non_bursting_master_requests <= internal_flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 OR internal_flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1;
  --pipeline_bridge_before_tristate_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pipeline_bridge_before_tristate_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pipeline_bridge_before_tristate_s1_arb_share_counter_next_value assignment, which is an e_assign
  pipeline_bridge_before_tristate_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pipeline_bridge_before_tristate_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_before_tristate_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(pipeline_bridge_before_tristate_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_before_tristate_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --pipeline_bridge_before_tristate_s1_allgrants all slave grants, which is an e_mux
  pipeline_bridge_before_tristate_s1_allgrants <= (pipeline_bridge_before_tristate_s1_grant_vector) OR (pipeline_bridge_before_tristate_s1_grant_vector);
  --pipeline_bridge_before_tristate_s1_end_xfer assignment, which is an e_assign
  pipeline_bridge_before_tristate_s1_end_xfer <= NOT ((pipeline_bridge_before_tristate_s1_waits_for_read OR pipeline_bridge_before_tristate_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_s1 <= pipeline_bridge_before_tristate_s1_end_xfer AND (((NOT pipeline_bridge_before_tristate_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pipeline_bridge_before_tristate_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pipeline_bridge_before_tristate_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_s1 AND pipeline_bridge_before_tristate_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_s1 AND NOT pipeline_bridge_before_tristate_s1_non_bursting_master_requests));
  --pipeline_bridge_before_tristate_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_before_tristate_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(pipeline_bridge_before_tristate_s1_arb_counter_enable) = '1' then 
        pipeline_bridge_before_tristate_s1_arb_share_counter <= pipeline_bridge_before_tristate_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pipeline_bridge_before_tristate_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_before_tristate_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pipeline_bridge_before_tristate_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_s1)) OR ((end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_s1 AND NOT pipeline_bridge_before_tristate_s1_non_bursting_master_requests)))) = '1' then 
        pipeline_bridge_before_tristate_s1_slavearbiterlockenable <= pipeline_bridge_before_tristate_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --flash_ssram_pipeline_bridge/m1 pipeline_bridge_before_tristate/s1 arbiterlock, which is an e_assign
  flash_ssram_pipeline_bridge_m1_arbiterlock <= pipeline_bridge_before_tristate_s1_slavearbiterlockenable AND flash_ssram_pipeline_bridge_m1_continuerequest;
  --pipeline_bridge_before_tristate_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pipeline_bridge_before_tristate_s1_slavearbiterlockenable2 <= pipeline_bridge_before_tristate_s1_arb_share_counter_next_value;
  --flash_ssram_pipeline_bridge/m1 pipeline_bridge_before_tristate/s1 arbiterlock2, which is an e_assign
  flash_ssram_pipeline_bridge_m1_arbiterlock2 <= pipeline_bridge_before_tristate_s1_slavearbiterlockenable2 AND flash_ssram_pipeline_bridge_m1_continuerequest;
  --pipeline_bridge_before_tristate_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pipeline_bridge_before_tristate_s1_any_continuerequest <= std_logic'('1');
  --flash_ssram_pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  flash_ssram_pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 <= internal_flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 AND NOT ((((flash_ssram_pipeline_bridge_m1_read AND flash_ssram_pipeline_bridge_m1_chipselect)) AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(flash_ssram_pipeline_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(flash_ssram_pipeline_bridge_m1_latency_counter))))))))));
  --unique name for pipeline_bridge_before_tristate_s1_move_on_to_next_transaction, which is an e_assign
  pipeline_bridge_before_tristate_s1_move_on_to_next_transaction <= pipeline_bridge_before_tristate_s1_readdatavalid_from_sa;
  --rdv_fifo_for_flash_ssram_pipeline_bridge_m1_to_pipeline_bridge_before_tristate_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_flash_ssram_pipeline_bridge_m1_to_pipeline_bridge_before_tristate_s1 : rdv_fifo_for_flash_ssram_pipeline_bridge_m1_to_pipeline_bridge_before_tristate_s1_module
    port map(
      data_out => flash_ssram_pipeline_bridge_m1_rdv_fifo_output_from_pipeline_bridge_before_tristate_s1,
      empty => open,
      fifo_contains_ones_n => flash_ssram_pipeline_bridge_m1_rdv_fifo_empty_pipeline_bridge_before_tristate_s1,
      full => open,
      clear_fifo => module_input22,
      clk => clk,
      data_in => internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1,
      read => pipeline_bridge_before_tristate_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input23,
      write => module_input24
    );

  module_input22 <= std_logic'('0');
  module_input23 <= std_logic'('0');
  module_input24 <= in_a_read_cycle AND NOT pipeline_bridge_before_tristate_s1_waits_for_read;

  flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1_shift_register <= NOT flash_ssram_pipeline_bridge_m1_rdv_fifo_empty_pipeline_bridge_before_tristate_s1;
  --local readdatavalid flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1, which is an e_mux
  flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1 <= pipeline_bridge_before_tristate_s1_readdatavalid_from_sa;
  --pipeline_bridge_before_tristate_s1_writedata mux, which is an e_mux
  pipeline_bridge_before_tristate_s1_writedata <= flash_ssram_pipeline_bridge_m1_writedata;
  --assign pipeline_bridge_before_tristate_s1_endofpacket_from_sa = pipeline_bridge_before_tristate_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  pipeline_bridge_before_tristate_s1_endofpacket_from_sa <= pipeline_bridge_before_tristate_s1_endofpacket;
  --master is always granted when requested
  internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 <= internal_flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1;
  --flash_ssram_pipeline_bridge/m1 saved-grant pipeline_bridge_before_tristate/s1, which is an e_assign
  flash_ssram_pipeline_bridge_m1_saved_grant_pipeline_bridge_before_tristate_s1 <= internal_flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1;
  --allow new arb cycle for pipeline_bridge_before_tristate/s1, which is an e_assign
  pipeline_bridge_before_tristate_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pipeline_bridge_before_tristate_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pipeline_bridge_before_tristate_s1_master_qreq_vector <= std_logic'('1');
  --pipeline_bridge_before_tristate_s1_reset_n assignment, which is an e_assign
  pipeline_bridge_before_tristate_s1_reset_n <= reset_n;
  pipeline_bridge_before_tristate_s1_chipselect <= internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1;
  --pipeline_bridge_before_tristate_s1_firsttransfer first transaction, which is an e_assign
  pipeline_bridge_before_tristate_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pipeline_bridge_before_tristate_s1_begins_xfer) = '1'), pipeline_bridge_before_tristate_s1_unreg_firsttransfer, pipeline_bridge_before_tristate_s1_reg_firsttransfer);
  --pipeline_bridge_before_tristate_s1_unreg_firsttransfer first transaction, which is an e_assign
  pipeline_bridge_before_tristate_s1_unreg_firsttransfer <= NOT ((pipeline_bridge_before_tristate_s1_slavearbiterlockenable AND pipeline_bridge_before_tristate_s1_any_continuerequest));
  --pipeline_bridge_before_tristate_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_before_tristate_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pipeline_bridge_before_tristate_s1_begins_xfer) = '1' then 
        pipeline_bridge_before_tristate_s1_reg_firsttransfer <= pipeline_bridge_before_tristate_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pipeline_bridge_before_tristate_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pipeline_bridge_before_tristate_s1_beginbursttransfer_internal <= pipeline_bridge_before_tristate_s1_begins_xfer;
  --pipeline_bridge_before_tristate_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  pipeline_bridge_before_tristate_s1_arbitration_holdoff_internal <= pipeline_bridge_before_tristate_s1_begins_xfer AND pipeline_bridge_before_tristate_s1_firsttransfer;
  --pipeline_bridge_before_tristate_s1_read assignment, which is an e_mux
  pipeline_bridge_before_tristate_s1_read <= internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 AND ((flash_ssram_pipeline_bridge_m1_read AND flash_ssram_pipeline_bridge_m1_chipselect));
  --pipeline_bridge_before_tristate_s1_write assignment, which is an e_mux
  pipeline_bridge_before_tristate_s1_write <= internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 AND ((flash_ssram_pipeline_bridge_m1_write AND flash_ssram_pipeline_bridge_m1_chipselect));
  shifted_address_to_pipeline_bridge_before_tristate_s1_from_flash_ssram_pipeline_bridge_m1 <= flash_ssram_pipeline_bridge_m1_address_to_slave;
  --pipeline_bridge_before_tristate_s1_address mux, which is an e_mux
  pipeline_bridge_before_tristate_s1_address <= A_EXT (A_SRL(shifted_address_to_pipeline_bridge_before_tristate_s1_from_flash_ssram_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 23);
  --slaveid pipeline_bridge_before_tristate_s1_nativeaddress nativeaddress mux, which is an e_mux
  pipeline_bridge_before_tristate_s1_nativeaddress <= A_EXT (A_SRL(flash_ssram_pipeline_bridge_m1_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 23);
  --d1_pipeline_bridge_before_tristate_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pipeline_bridge_before_tristate_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pipeline_bridge_before_tristate_s1_end_xfer <= pipeline_bridge_before_tristate_s1_end_xfer;
    end if;

  end process;

  --pipeline_bridge_before_tristate_s1_waits_for_read in a cycle, which is an e_mux
  pipeline_bridge_before_tristate_s1_waits_for_read <= pipeline_bridge_before_tristate_s1_in_a_read_cycle AND internal_pipeline_bridge_before_tristate_s1_waitrequest_from_sa;
  --pipeline_bridge_before_tristate_s1_in_a_read_cycle assignment, which is an e_assign
  pipeline_bridge_before_tristate_s1_in_a_read_cycle <= internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 AND ((flash_ssram_pipeline_bridge_m1_read AND flash_ssram_pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pipeline_bridge_before_tristate_s1_in_a_read_cycle;
  --pipeline_bridge_before_tristate_s1_waits_for_write in a cycle, which is an e_mux
  pipeline_bridge_before_tristate_s1_waits_for_write <= pipeline_bridge_before_tristate_s1_in_a_write_cycle AND internal_pipeline_bridge_before_tristate_s1_waitrequest_from_sa;
  --pipeline_bridge_before_tristate_s1_in_a_write_cycle assignment, which is an e_assign
  pipeline_bridge_before_tristate_s1_in_a_write_cycle <= internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 AND ((flash_ssram_pipeline_bridge_m1_write AND flash_ssram_pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pipeline_bridge_before_tristate_s1_in_a_write_cycle;
  wait_for_pipeline_bridge_before_tristate_s1_counter <= std_logic'('0');
  --pipeline_bridge_before_tristate_s1_byteenable byte enable port mux, which is an e_mux
  pipeline_bridge_before_tristate_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (flash_ssram_pipeline_bridge_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  pipeline_bridge_before_tristate_s1_burstcount <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(flash_ssram_pipeline_bridge_m1_burstcount))), std_logic_vector'("00000000000000000000000000000001")));
  --pipeline_bridge_before_tristate/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  pipeline_bridge_before_tristate_s1_arbiterlock <= flash_ssram_pipeline_bridge_m1_arbiterlock;
  --pipeline_bridge_before_tristate/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  pipeline_bridge_before_tristate_s1_arbiterlock2 <= flash_ssram_pipeline_bridge_m1_arbiterlock2;
  --debugaccess mux, which is an e_mux
  pipeline_bridge_before_tristate_s1_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(flash_ssram_pipeline_bridge_m1_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 <= internal_flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1;
  --vhdl renameroo for output signals
  flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 <= internal_flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1;
  --vhdl renameroo for output signals
  flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 <= internal_flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_s1_waitrequest_from_sa <= internal_pipeline_bridge_before_tristate_s1_waitrequest_from_sa;
--synthesis translate_off
    --pipeline_bridge_before_tristate/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --flash_ssram_pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line52 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(flash_ssram_pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line52, now);
          write(write_line52, string'(": "));
          write(write_line52, string'("flash_ssram_pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave pipeline_bridge_before_tristate/s1"));
          write(output, write_line52.all);
          deallocate (write_line52);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pipeline_bridge_before_tristate_m1_arbitrator is 
        port (
              -- inputs:
                 signal cfi_flash_s1_wait_counter_eq_0 : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal d1_flash_ssram_tristate_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal incoming_flash_ssram_tristate_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal incoming_flash_ssram_tristate_data_with_Xs_converted_to_0 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_granted_ssram_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_requests_ssram_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal pipeline_bridge_before_tristate_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_latency_counter : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_before_tristate_m1_readdatavalid : OUT STD_LOGIC;
                 signal pipeline_bridge_before_tristate_m1_waitrequest : OUT STD_LOGIC
              );
end entity pipeline_bridge_before_tristate_m1_arbitrator;


architecture europa of pipeline_bridge_before_tristate_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_pipeline_bridge_before_tristate_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_pipeline_bridge_before_tristate_m1_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_pipeline_bridge_before_tristate_m1_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_pipeline_bridge_before_tristate_m1_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_pipeline_bridge_before_tristate_m1_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_burstcount_last_time :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_chipselect_last_time :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_is_granted_some_slave :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_read_but_no_slave_selected :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_read_last_time :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_run :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_write_last_time :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_pipeline_bridge_before_tristate_m1_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 OR (((((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect)) AND NOT(or_reduce(pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1))) AND internal_pipeline_bridge_before_tristate_m1_dbs_address(1)))) OR NOT pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 OR NOT pipeline_bridge_before_tristate_m1_requests_ssram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 OR NOT ((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect)))))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cfi_flash_s1_wait_counter_eq_0 AND NOT d1_flash_ssram_tristate_avalon_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_pipeline_bridge_before_tristate_m1_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 OR NOT ((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect)))))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cfi_flash_s1_wait_counter_eq_0 AND NOT d1_flash_ssram_tristate_avalon_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_pipeline_bridge_before_tristate_m1_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 OR NOT pipeline_bridge_before_tristate_m1_chipselect)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_before_tristate_m1_chipselect)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 OR NOT pipeline_bridge_before_tristate_m1_chipselect)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_before_tristate_m1_chipselect)))))))));
  --cascaded wait assignment, which is an e_assign
  pipeline_bridge_before_tristate_m1_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_pipeline_bridge_before_tristate_m1_address_to_slave <= pipeline_bridge_before_tristate_m1_address(24 DOWNTO 0);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic((((((((NOT std_logic_vector'("00000000000000000000000000000000")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT(or_reduce(pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1))))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 AND ((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect)))))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cfi_flash_s1_wait_counter_eq_0 AND NOT d1_flash_ssram_tristate_avalon_slave_end_xfer)))))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 AND ((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect)))))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cfi_flash_s1_wait_counter_eq_0 AND NOT d1_flash_ssram_tristate_avalon_slave_end_xfer)))))))));
  --pipeline_bridge_before_tristate_m1_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_before_tristate_m1_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pipeline_bridge_before_tristate_m1_read_but_no_slave_selected <= (((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect)) AND pipeline_bridge_before_tristate_m1_run) AND NOT pipeline_bridge_before_tristate_m1_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  pipeline_bridge_before_tristate_m1_is_granted_some_slave <= pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 OR pipeline_bridge_before_tristate_m1_granted_ssram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pipeline_bridge_before_tristate_m1_readdatavalid <= ((pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1 AND dbs_rdv_counter_overflow)) OR pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  pipeline_bridge_before_tristate_m1_readdatavalid <= ((pipeline_bridge_before_tristate_m1_read_but_no_slave_selected OR pre_flush_pipeline_bridge_before_tristate_m1_readdatavalid) OR pipeline_bridge_before_tristate_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_before_tristate_m1_readdatavalid;
  --input to latent dbs-16 stored 0, which is an e_mux
  p1_dbs_latent_16_reg_segment_0 <= incoming_flash_ssram_tristate_data_with_Xs_converted_to_0;
  --dbs register for latent dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pipeline_bridge_before_tristate_m1_dbs_rdv_counter(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
      end if;
    end if;

  end process;

  --pipeline_bridge_before_tristate/m1 readdata mux, which is an e_mux
  pipeline_bridge_before_tristate_m1_readdata <= ((A_REP(NOT pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1, 32) OR Std_Logic_Vector'(incoming_flash_ssram_tristate_data_with_Xs_converted_to_0(15 DOWNTO 0) & dbs_latent_16_reg_segment_0))) AND ((A_REP(NOT pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1, 32) OR incoming_flash_ssram_tristate_data));
  --mux write dbs 1, which is an e_mux
  pipeline_bridge_before_tristate_m1_dbs_write_16 <= A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_before_tristate_m1_dbs_address(1))) = '1'), pipeline_bridge_before_tristate_m1_writedata(31 DOWNTO 16), pipeline_bridge_before_tristate_m1_writedata(15 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_pipeline_bridge_before_tristate_m1_waitrequest <= NOT pipeline_bridge_before_tristate_m1_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pipeline_bridge_before_tristate_m1_latency_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      internal_pipeline_bridge_before_tristate_m1_latency_counter <= p1_pipeline_bridge_before_tristate_m1_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_pipeline_bridge_before_tristate_m1_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((pipeline_bridge_before_tristate_m1_run AND ((pipeline_bridge_before_tristate_m1_read AND pipeline_bridge_before_tristate_m1_chipselect))))) = '1'), (std_logic_vector'("000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_pipeline_bridge_before_tristate_m1_latency_counter)) /= std_logic_vector'("000")), ((std_logic_vector'("000000000000000000000000000000") & (internal_pipeline_bridge_before_tristate_m1_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT (((((std_logic_vector'("00000000000000000000000000000") & (A_REP(pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1, 3))) AND std_logic_vector'("00000000000000000000000000000010"))) OR (((std_logic_vector'("00000000000000000000000000000") & (A_REP(pipeline_bridge_before_tristate_m1_requests_ssram_s1, 3))) AND std_logic_vector'("00000000000000000000000000000100")))), 3);
  --dbs count increment, which is an e_mux
  pipeline_bridge_before_tristate_m1_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_pipeline_bridge_before_tristate_m1_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_pipeline_bridge_before_tristate_m1_dbs_address)) + (std_logic_vector'("0") & (pipeline_bridge_before_tristate_m1_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pipeline_bridge_before_tristate_m1_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_pipeline_bridge_before_tristate_m1_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  pipeline_bridge_before_tristate_m1_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (pipeline_bridge_before_tristate_m1_dbs_rdv_counter)) + (std_logic_vector'("0") & (pipeline_bridge_before_tristate_m1_dbs_rdv_counter_inc))), 2);
  --pipeline_bridge_before_tristate_m1_rdv_inc_mux, which is an e_mux
  pipeline_bridge_before_tristate_m1_dbs_rdv_counter_inc <= std_logic_vector'("10");
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_before_tristate_m1_dbs_rdv_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        pipeline_bridge_before_tristate_m1_dbs_rdv_counter <= pipeline_bridge_before_tristate_m1_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= pipeline_bridge_before_tristate_m1_dbs_rdv_counter(1) AND NOT pipeline_bridge_before_tristate_m1_next_dbs_rdv_counter(1);
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_address_to_slave <= internal_pipeline_bridge_before_tristate_m1_address_to_slave;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_dbs_address <= internal_pipeline_bridge_before_tristate_m1_dbs_address;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_latency_counter <= internal_pipeline_bridge_before_tristate_m1_latency_counter;
  --vhdl renameroo for output signals
  pipeline_bridge_before_tristate_m1_waitrequest <= internal_pipeline_bridge_before_tristate_m1_waitrequest;
--synthesis translate_off
    --pipeline_bridge_before_tristate_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_before_tristate_m1_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        pipeline_bridge_before_tristate_m1_address_last_time <= pipeline_bridge_before_tristate_m1_address;
      end if;

    end process;

    --pipeline_bridge_before_tristate/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pipeline_bridge_before_tristate_m1_waitrequest AND pipeline_bridge_before_tristate_m1_chipselect;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line53 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pipeline_bridge_before_tristate_m1_address /= pipeline_bridge_before_tristate_m1_address_last_time))))) = '1' then 
          write(write_line53, now);
          write(write_line53, string'(": "));
          write(write_line53, string'("pipeline_bridge_before_tristate_m1_address did not heed wait!!!"));
          write(output, write_line53.all);
          deallocate (write_line53);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_chipselect check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_before_tristate_m1_chipselect_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pipeline_bridge_before_tristate_m1_chipselect_last_time <= pipeline_bridge_before_tristate_m1_chipselect;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_chipselect matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line54 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pipeline_bridge_before_tristate_m1_chipselect) /= std_logic'(pipeline_bridge_before_tristate_m1_chipselect_last_time)))))) = '1' then 
          write(write_line54, now);
          write(write_line54, string'(": "));
          write(write_line54, string'("pipeline_bridge_before_tristate_m1_chipselect did not heed wait!!!"));
          write(output, write_line54.all);
          deallocate (write_line54);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_before_tristate_m1_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pipeline_bridge_before_tristate_m1_burstcount_last_time <= pipeline_bridge_before_tristate_m1_burstcount;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line55 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pipeline_bridge_before_tristate_m1_burstcount) /= std_logic'(pipeline_bridge_before_tristate_m1_burstcount_last_time)))))) = '1' then 
          write(write_line55, now);
          write(write_line55, string'(": "));
          write(write_line55, string'("pipeline_bridge_before_tristate_m1_burstcount did not heed wait!!!"));
          write(output, write_line55.all);
          deallocate (write_line55);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_before_tristate_m1_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        pipeline_bridge_before_tristate_m1_byteenable_last_time <= pipeline_bridge_before_tristate_m1_byteenable;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line56 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pipeline_bridge_before_tristate_m1_byteenable /= pipeline_bridge_before_tristate_m1_byteenable_last_time))))) = '1' then 
          write(write_line56, now);
          write(write_line56, string'(": "));
          write(write_line56, string'("pipeline_bridge_before_tristate_m1_byteenable did not heed wait!!!"));
          write(output, write_line56.all);
          deallocate (write_line56);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_before_tristate_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pipeline_bridge_before_tristate_m1_read_last_time <= pipeline_bridge_before_tristate_m1_read;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line57 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pipeline_bridge_before_tristate_m1_read) /= std_logic'(pipeline_bridge_before_tristate_m1_read_last_time)))))) = '1' then 
          write(write_line57, now);
          write(write_line57, string'(": "));
          write(write_line57, string'("pipeline_bridge_before_tristate_m1_read did not heed wait!!!"));
          write(output, write_line57.all);
          deallocate (write_line57);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_before_tristate_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pipeline_bridge_before_tristate_m1_write_last_time <= pipeline_bridge_before_tristate_m1_write;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line58 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pipeline_bridge_before_tristate_m1_write) /= std_logic'(pipeline_bridge_before_tristate_m1_write_last_time)))))) = '1' then 
          write(write_line58, now);
          write(write_line58, string'(": "));
          write(write_line58, string'("pipeline_bridge_before_tristate_m1_write did not heed wait!!!"));
          write(output, write_line58.all);
          deallocate (write_line58);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_before_tristate_m1_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pipeline_bridge_before_tristate_m1_writedata_last_time <= pipeline_bridge_before_tristate_m1_writedata;
      end if;

    end process;

    --pipeline_bridge_before_tristate_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line59 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((pipeline_bridge_before_tristate_m1_writedata /= pipeline_bridge_before_tristate_m1_writedata_last_time)))) AND ((pipeline_bridge_before_tristate_m1_write AND pipeline_bridge_before_tristate_m1_chipselect)))) = '1' then 
          write(write_line59, now);
          write(write_line59, string'(": "));
          write(write_line59, string'("pipeline_bridge_before_tristate_m1_writedata did not heed wait!!!"));
          write(output, write_line59.all);
          deallocate (write_line59);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pipeline_bridge_before_tristate_bridge_arbitrator is 
end entity pipeline_bridge_before_tristate_bridge_arbitrator;


architecture europa of pipeline_bridge_before_tristate_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pll_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal gpib_edm1_clock_0_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal gpib_edm1_clock_0_out_read : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_out_write : IN STD_LOGIC;
                 signal gpib_edm1_clock_0_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pll_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pll_s1_resetrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pll_s1_end_xfer : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_out_granted_pll_s1 : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_out_qualified_request_pll_s1 : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_out_read_data_valid_pll_s1 : OUT STD_LOGIC;
                 signal gpib_edm1_clock_0_out_requests_pll_s1 : OUT STD_LOGIC;
                 signal pll_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal pll_s1_chipselect : OUT STD_LOGIC;
                 signal pll_s1_read : OUT STD_LOGIC;
                 signal pll_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pll_s1_reset_n : OUT STD_LOGIC;
                 signal pll_s1_resetrequest_from_sa : OUT STD_LOGIC;
                 signal pll_s1_write : OUT STD_LOGIC;
                 signal pll_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pll_s1_arbitrator;


architecture europa of pll_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pll_s1 :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_arbiterlock :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_arbiterlock2 :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_continuerequest :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_saved_grant_pll_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_gpib_edm1_clock_0_out_granted_pll_s1 :  STD_LOGIC;
                signal internal_gpib_edm1_clock_0_out_qualified_request_pll_s1 :  STD_LOGIC;
                signal internal_gpib_edm1_clock_0_out_requests_pll_s1 :  STD_LOGIC;
                signal pll_s1_allgrants :  STD_LOGIC;
                signal pll_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pll_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pll_s1_any_continuerequest :  STD_LOGIC;
                signal pll_s1_arb_counter_enable :  STD_LOGIC;
                signal pll_s1_arb_share_counter :  STD_LOGIC;
                signal pll_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal pll_s1_arb_share_set_values :  STD_LOGIC;
                signal pll_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pll_s1_begins_xfer :  STD_LOGIC;
                signal pll_s1_end_xfer :  STD_LOGIC;
                signal pll_s1_firsttransfer :  STD_LOGIC;
                signal pll_s1_grant_vector :  STD_LOGIC;
                signal pll_s1_in_a_read_cycle :  STD_LOGIC;
                signal pll_s1_in_a_write_cycle :  STD_LOGIC;
                signal pll_s1_master_qreq_vector :  STD_LOGIC;
                signal pll_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pll_s1_reg_firsttransfer :  STD_LOGIC;
                signal pll_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pll_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pll_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pll_s1_waits_for_read :  STD_LOGIC;
                signal pll_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_pll_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pll_s1_end_xfer;
    end if;

  end process;

  pll_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_gpib_edm1_clock_0_out_qualified_request_pll_s1);
  --assign pll_s1_readdata_from_sa = pll_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pll_s1_readdata_from_sa <= pll_s1_readdata;
  internal_gpib_edm1_clock_0_out_requests_pll_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((gpib_edm1_clock_0_out_read OR gpib_edm1_clock_0_out_write)))))));
  --pll_s1_arb_share_counter set values, which is an e_mux
  pll_s1_arb_share_set_values <= std_logic'('1');
  --pll_s1_non_bursting_master_requests mux, which is an e_mux
  pll_s1_non_bursting_master_requests <= internal_gpib_edm1_clock_0_out_requests_pll_s1;
  --pll_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pll_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pll_s1_arb_share_counter_next_value assignment, which is an e_assign
  pll_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pll_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pll_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(pll_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pll_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --pll_s1_allgrants all slave grants, which is an e_mux
  pll_s1_allgrants <= pll_s1_grant_vector;
  --pll_s1_end_xfer assignment, which is an e_assign
  pll_s1_end_xfer <= NOT ((pll_s1_waits_for_read OR pll_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pll_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pll_s1 <= pll_s1_end_xfer AND (((NOT pll_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pll_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pll_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pll_s1 AND pll_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pll_s1 AND NOT pll_s1_non_bursting_master_requests));
  --pll_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pll_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(pll_s1_arb_counter_enable) = '1' then 
        pll_s1_arb_share_counter <= pll_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pll_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pll_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pll_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pll_s1)) OR ((end_xfer_arb_share_counter_term_pll_s1 AND NOT pll_s1_non_bursting_master_requests)))) = '1' then 
        pll_s1_slavearbiterlockenable <= pll_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_0/out pll/s1 arbiterlock, which is an e_assign
  gpib_edm1_clock_0_out_arbiterlock <= pll_s1_slavearbiterlockenable AND gpib_edm1_clock_0_out_continuerequest;
  --pll_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pll_s1_slavearbiterlockenable2 <= pll_s1_arb_share_counter_next_value;
  --gpib_edm1_clock_0/out pll/s1 arbiterlock2, which is an e_assign
  gpib_edm1_clock_0_out_arbiterlock2 <= pll_s1_slavearbiterlockenable2 AND gpib_edm1_clock_0_out_continuerequest;
  --pll_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pll_s1_any_continuerequest <= std_logic'('1');
  --gpib_edm1_clock_0_out_continuerequest continued request, which is an e_assign
  gpib_edm1_clock_0_out_continuerequest <= std_logic'('1');
  internal_gpib_edm1_clock_0_out_qualified_request_pll_s1 <= internal_gpib_edm1_clock_0_out_requests_pll_s1;
  --pll_s1_writedata mux, which is an e_mux
  pll_s1_writedata <= gpib_edm1_clock_0_out_writedata;
  --master is always granted when requested
  internal_gpib_edm1_clock_0_out_granted_pll_s1 <= internal_gpib_edm1_clock_0_out_qualified_request_pll_s1;
  --gpib_edm1_clock_0/out saved-grant pll/s1, which is an e_assign
  gpib_edm1_clock_0_out_saved_grant_pll_s1 <= internal_gpib_edm1_clock_0_out_requests_pll_s1;
  --allow new arb cycle for pll/s1, which is an e_assign
  pll_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pll_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pll_s1_master_qreq_vector <= std_logic'('1');
  --pll_s1_reset_n assignment, which is an e_assign
  pll_s1_reset_n <= reset_n;
  --assign pll_s1_resetrequest_from_sa = pll_s1_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  pll_s1_resetrequest_from_sa <= pll_s1_resetrequest;
  pll_s1_chipselect <= internal_gpib_edm1_clock_0_out_granted_pll_s1;
  --pll_s1_firsttransfer first transaction, which is an e_assign
  pll_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pll_s1_begins_xfer) = '1'), pll_s1_unreg_firsttransfer, pll_s1_reg_firsttransfer);
  --pll_s1_unreg_firsttransfer first transaction, which is an e_assign
  pll_s1_unreg_firsttransfer <= NOT ((pll_s1_slavearbiterlockenable AND pll_s1_any_continuerequest));
  --pll_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pll_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pll_s1_begins_xfer) = '1' then 
        pll_s1_reg_firsttransfer <= pll_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pll_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pll_s1_beginbursttransfer_internal <= pll_s1_begins_xfer;
  --pll_s1_read assignment, which is an e_mux
  pll_s1_read <= internal_gpib_edm1_clock_0_out_granted_pll_s1 AND gpib_edm1_clock_0_out_read;
  --pll_s1_write assignment, which is an e_mux
  pll_s1_write <= internal_gpib_edm1_clock_0_out_granted_pll_s1 AND gpib_edm1_clock_0_out_write;
  --pll_s1_address mux, which is an e_mux
  pll_s1_address <= gpib_edm1_clock_0_out_nativeaddress;
  --d1_pll_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pll_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pll_s1_end_xfer <= pll_s1_end_xfer;
    end if;

  end process;

  --pll_s1_waits_for_read in a cycle, which is an e_mux
  pll_s1_waits_for_read <= pll_s1_in_a_read_cycle AND pll_s1_begins_xfer;
  --pll_s1_in_a_read_cycle assignment, which is an e_assign
  pll_s1_in_a_read_cycle <= internal_gpib_edm1_clock_0_out_granted_pll_s1 AND gpib_edm1_clock_0_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pll_s1_in_a_read_cycle;
  --pll_s1_waits_for_write in a cycle, which is an e_mux
  pll_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pll_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pll_s1_in_a_write_cycle assignment, which is an e_assign
  pll_s1_in_a_write_cycle <= internal_gpib_edm1_clock_0_out_granted_pll_s1 AND gpib_edm1_clock_0_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pll_s1_in_a_write_cycle;
  wait_for_pll_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  gpib_edm1_clock_0_out_granted_pll_s1 <= internal_gpib_edm1_clock_0_out_granted_pll_s1;
  --vhdl renameroo for output signals
  gpib_edm1_clock_0_out_qualified_request_pll_s1 <= internal_gpib_edm1_clock_0_out_qualified_request_pll_s1;
  --vhdl renameroo for output signals
  gpib_edm1_clock_0_out_requests_pll_s1 <= internal_gpib_edm1_clock_0_out_requests_pll_s1;
--synthesis translate_off
    --pll/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity remote_update_cycloneiii_1_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_out_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gpib_edm1_clock_1_out_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal gpib_edm1_clock_1_out_read : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_out_write : IN STD_LOGIC;
                 signal gpib_edm1_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal remote_update_cycloneiii_1_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal remote_update_cycloneiii_1_s1_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_remote_update_cycloneiii_1_s1_end_xfer : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1 : OUT STD_LOGIC;
                 signal gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_1_s1_address : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal remote_update_cycloneiii_1_s1_chipselect : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_1_s1_read : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal remote_update_cycloneiii_1_s1_reset : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_1_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_1_s1_write : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_1_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity remote_update_cycloneiii_1_s1_arbitrator;


architecture europa of remote_update_cycloneiii_1_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_remote_update_cycloneiii_1_s1 :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_arbiterlock :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_arbiterlock2 :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_continuerequest :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register_in :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_saved_grant_remote_update_cycloneiii_1_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 :  STD_LOGIC;
                signal internal_gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 :  STD_LOGIC;
                signal internal_gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 :  STD_LOGIC;
                signal internal_remote_update_cycloneiii_1_s1_waitrequest_from_sa :  STD_LOGIC;
                signal p1_gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal remote_update_cycloneiii_1_s1_allgrants :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_any_continuerequest :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_arb_counter_enable :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_arb_share_counter :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_arb_share_set_values :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_begins_xfer :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_end_xfer :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_firsttransfer :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_grant_vector :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_in_a_read_cycle :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_in_a_write_cycle :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_master_qreq_vector :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_non_bursting_master_requests :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_reg_firsttransfer :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_slavearbiterlockenable :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_unreg_firsttransfer :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_waits_for_read :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_remote_update_cycloneiii_1_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT remote_update_cycloneiii_1_s1_end_xfer;
    end if;

  end process;

  remote_update_cycloneiii_1_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1);
  --assign remote_update_cycloneiii_1_s1_readdata_from_sa = remote_update_cycloneiii_1_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  remote_update_cycloneiii_1_s1_readdata_from_sa <= remote_update_cycloneiii_1_s1_readdata;
  internal_gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((gpib_edm1_clock_1_out_read OR gpib_edm1_clock_1_out_write)))))));
  --assign remote_update_cycloneiii_1_s1_waitrequest_from_sa = remote_update_cycloneiii_1_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_remote_update_cycloneiii_1_s1_waitrequest_from_sa <= remote_update_cycloneiii_1_s1_waitrequest;
  --remote_update_cycloneiii_1_s1_arb_share_counter set values, which is an e_mux
  remote_update_cycloneiii_1_s1_arb_share_set_values <= std_logic'('1');
  --remote_update_cycloneiii_1_s1_non_bursting_master_requests mux, which is an e_mux
  remote_update_cycloneiii_1_s1_non_bursting_master_requests <= internal_gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1;
  --remote_update_cycloneiii_1_s1_any_bursting_master_saved_grant mux, which is an e_mux
  remote_update_cycloneiii_1_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --remote_update_cycloneiii_1_s1_arb_share_counter_next_value assignment, which is an e_assign
  remote_update_cycloneiii_1_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(remote_update_cycloneiii_1_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(remote_update_cycloneiii_1_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(remote_update_cycloneiii_1_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(remote_update_cycloneiii_1_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --remote_update_cycloneiii_1_s1_allgrants all slave grants, which is an e_mux
  remote_update_cycloneiii_1_s1_allgrants <= remote_update_cycloneiii_1_s1_grant_vector;
  --remote_update_cycloneiii_1_s1_end_xfer assignment, which is an e_assign
  remote_update_cycloneiii_1_s1_end_xfer <= NOT ((remote_update_cycloneiii_1_s1_waits_for_read OR remote_update_cycloneiii_1_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_remote_update_cycloneiii_1_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_remote_update_cycloneiii_1_s1 <= remote_update_cycloneiii_1_s1_end_xfer AND (((NOT remote_update_cycloneiii_1_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --remote_update_cycloneiii_1_s1_arb_share_counter arbitration counter enable, which is an e_assign
  remote_update_cycloneiii_1_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_remote_update_cycloneiii_1_s1 AND remote_update_cycloneiii_1_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_remote_update_cycloneiii_1_s1 AND NOT remote_update_cycloneiii_1_s1_non_bursting_master_requests));
  --remote_update_cycloneiii_1_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      remote_update_cycloneiii_1_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(remote_update_cycloneiii_1_s1_arb_counter_enable) = '1' then 
        remote_update_cycloneiii_1_s1_arb_share_counter <= remote_update_cycloneiii_1_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --remote_update_cycloneiii_1_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      remote_update_cycloneiii_1_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((remote_update_cycloneiii_1_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_remote_update_cycloneiii_1_s1)) OR ((end_xfer_arb_share_counter_term_remote_update_cycloneiii_1_s1 AND NOT remote_update_cycloneiii_1_s1_non_bursting_master_requests)))) = '1' then 
        remote_update_cycloneiii_1_s1_slavearbiterlockenable <= remote_update_cycloneiii_1_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --gpib_edm1_clock_1/out remote_update_cycloneiii_1/s1 arbiterlock, which is an e_assign
  gpib_edm1_clock_1_out_arbiterlock <= remote_update_cycloneiii_1_s1_slavearbiterlockenable AND gpib_edm1_clock_1_out_continuerequest;
  --remote_update_cycloneiii_1_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  remote_update_cycloneiii_1_s1_slavearbiterlockenable2 <= remote_update_cycloneiii_1_s1_arb_share_counter_next_value;
  --gpib_edm1_clock_1/out remote_update_cycloneiii_1/s1 arbiterlock2, which is an e_assign
  gpib_edm1_clock_1_out_arbiterlock2 <= remote_update_cycloneiii_1_s1_slavearbiterlockenable2 AND gpib_edm1_clock_1_out_continuerequest;
  --remote_update_cycloneiii_1_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  remote_update_cycloneiii_1_s1_any_continuerequest <= std_logic'('1');
  --gpib_edm1_clock_1_out_continuerequest continued request, which is an e_assign
  gpib_edm1_clock_1_out_continuerequest <= std_logic'('1');
  internal_gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 <= internal_gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 AND NOT ((gpib_edm1_clock_1_out_read AND (or_reduce(gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register))));
  --gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register_in <= ((internal_gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 AND gpib_edm1_clock_1_out_read) AND NOT remote_update_cycloneiii_1_s1_waits_for_read) AND NOT (or_reduce(gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register));
  --shift register p1 gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register <= A_EXT ((gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register & A_ToStdLogicVector(gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register_in)), 2);
  --gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register <= p1_gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register;
    end if;

  end process;

  --local readdatavalid gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1, which is an e_mux
  gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1 <= gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1_shift_register(1);
  --remote_update_cycloneiii_1_s1_writedata mux, which is an e_mux
  remote_update_cycloneiii_1_s1_writedata <= gpib_edm1_clock_1_out_writedata;
  --master is always granted when requested
  internal_gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 <= internal_gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1;
  --gpib_edm1_clock_1/out saved-grant remote_update_cycloneiii_1/s1, which is an e_assign
  gpib_edm1_clock_1_out_saved_grant_remote_update_cycloneiii_1_s1 <= internal_gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1;
  --allow new arb cycle for remote_update_cycloneiii_1/s1, which is an e_assign
  remote_update_cycloneiii_1_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  remote_update_cycloneiii_1_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  remote_update_cycloneiii_1_s1_master_qreq_vector <= std_logic'('1');
  --~remote_update_cycloneiii_1_s1_reset assignment, which is an e_assign
  remote_update_cycloneiii_1_s1_reset <= NOT reset_n;
  remote_update_cycloneiii_1_s1_chipselect <= internal_gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1;
  --remote_update_cycloneiii_1_s1_firsttransfer first transaction, which is an e_assign
  remote_update_cycloneiii_1_s1_firsttransfer <= A_WE_StdLogic((std_logic'(remote_update_cycloneiii_1_s1_begins_xfer) = '1'), remote_update_cycloneiii_1_s1_unreg_firsttransfer, remote_update_cycloneiii_1_s1_reg_firsttransfer);
  --remote_update_cycloneiii_1_s1_unreg_firsttransfer first transaction, which is an e_assign
  remote_update_cycloneiii_1_s1_unreg_firsttransfer <= NOT ((remote_update_cycloneiii_1_s1_slavearbiterlockenable AND remote_update_cycloneiii_1_s1_any_continuerequest));
  --remote_update_cycloneiii_1_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      remote_update_cycloneiii_1_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(remote_update_cycloneiii_1_s1_begins_xfer) = '1' then 
        remote_update_cycloneiii_1_s1_reg_firsttransfer <= remote_update_cycloneiii_1_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --remote_update_cycloneiii_1_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  remote_update_cycloneiii_1_s1_beginbursttransfer_internal <= remote_update_cycloneiii_1_s1_begins_xfer;
  --remote_update_cycloneiii_1_s1_read assignment, which is an e_mux
  remote_update_cycloneiii_1_s1_read <= internal_gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 AND gpib_edm1_clock_1_out_read;
  --remote_update_cycloneiii_1_s1_write assignment, which is an e_mux
  remote_update_cycloneiii_1_s1_write <= internal_gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 AND gpib_edm1_clock_1_out_write;
  --remote_update_cycloneiii_1_s1_address mux, which is an e_mux
  remote_update_cycloneiii_1_s1_address <= gpib_edm1_clock_1_out_nativeaddress;
  --d1_remote_update_cycloneiii_1_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_remote_update_cycloneiii_1_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_remote_update_cycloneiii_1_s1_end_xfer <= remote_update_cycloneiii_1_s1_end_xfer;
    end if;

  end process;

  --remote_update_cycloneiii_1_s1_waits_for_read in a cycle, which is an e_mux
  remote_update_cycloneiii_1_s1_waits_for_read <= remote_update_cycloneiii_1_s1_in_a_read_cycle AND internal_remote_update_cycloneiii_1_s1_waitrequest_from_sa;
  --remote_update_cycloneiii_1_s1_in_a_read_cycle assignment, which is an e_assign
  remote_update_cycloneiii_1_s1_in_a_read_cycle <= internal_gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 AND gpib_edm1_clock_1_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= remote_update_cycloneiii_1_s1_in_a_read_cycle;
  --remote_update_cycloneiii_1_s1_waits_for_write in a cycle, which is an e_mux
  remote_update_cycloneiii_1_s1_waits_for_write <= remote_update_cycloneiii_1_s1_in_a_write_cycle AND internal_remote_update_cycloneiii_1_s1_waitrequest_from_sa;
  --remote_update_cycloneiii_1_s1_in_a_write_cycle assignment, which is an e_assign
  remote_update_cycloneiii_1_s1_in_a_write_cycle <= internal_gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 AND gpib_edm1_clock_1_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= remote_update_cycloneiii_1_s1_in_a_write_cycle;
  wait_for_remote_update_cycloneiii_1_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 <= internal_gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1;
  --vhdl renameroo for output signals
  gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 <= internal_gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1;
  --vhdl renameroo for output signals
  gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 <= internal_gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1;
  --vhdl renameroo for output signals
  remote_update_cycloneiii_1_s1_waitrequest_from_sa <= internal_remote_update_cycloneiii_1_s1_waitrequest_from_sa;
--synthesis translate_off
    --remote_update_cycloneiii_1/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sys_clk_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_s1_irq : IN STD_LOGIC;
                 signal sys_clk_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal clock_crossing_0_m1_granted_sys_clk_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_sys_clk_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_sys_clk_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_sys_clk_s1 : OUT STD_LOGIC;
                 signal d1_sys_clk_s1_end_xfer : OUT STD_LOGIC;
                 signal sys_clk_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal sys_clk_s1_chipselect : OUT STD_LOGIC;
                 signal sys_clk_s1_irq_from_sa : OUT STD_LOGIC;
                 signal sys_clk_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sys_clk_s1_reset_n : OUT STD_LOGIC;
                 signal sys_clk_s1_write_n : OUT STD_LOGIC;
                 signal sys_clk_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sys_clk_s1_arbitrator;


architecture europa of sys_clk_s1_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_sys_clk_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sys_clk_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_sys_clk_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_sys_clk_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_sys_clk_s1 :  STD_LOGIC;
                signal sys_clk_s1_allgrants :  STD_LOGIC;
                signal sys_clk_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sys_clk_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sys_clk_s1_any_continuerequest :  STD_LOGIC;
                signal sys_clk_s1_arb_counter_enable :  STD_LOGIC;
                signal sys_clk_s1_arb_share_counter :  STD_LOGIC;
                signal sys_clk_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal sys_clk_s1_arb_share_set_values :  STD_LOGIC;
                signal sys_clk_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sys_clk_s1_begins_xfer :  STD_LOGIC;
                signal sys_clk_s1_end_xfer :  STD_LOGIC;
                signal sys_clk_s1_firsttransfer :  STD_LOGIC;
                signal sys_clk_s1_grant_vector :  STD_LOGIC;
                signal sys_clk_s1_in_a_read_cycle :  STD_LOGIC;
                signal sys_clk_s1_in_a_write_cycle :  STD_LOGIC;
                signal sys_clk_s1_master_qreq_vector :  STD_LOGIC;
                signal sys_clk_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sys_clk_s1_reg_firsttransfer :  STD_LOGIC;
                signal sys_clk_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sys_clk_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sys_clk_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sys_clk_s1_waits_for_read :  STD_LOGIC;
                signal sys_clk_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_sys_clk_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sys_clk_s1_end_xfer;
    end if;

  end process;

  sys_clk_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_sys_clk_s1);
  --assign sys_clk_s1_readdata_from_sa = sys_clk_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sys_clk_s1_readdata_from_sa <= sys_clk_s1_readdata;
  internal_clock_crossing_0_m1_requests_sys_clk_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(7 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("00000000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --sys_clk_s1_arb_share_counter set values, which is an e_mux
  sys_clk_s1_arb_share_set_values <= std_logic'('1');
  --sys_clk_s1_non_bursting_master_requests mux, which is an e_mux
  sys_clk_s1_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_sys_clk_s1;
  --sys_clk_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sys_clk_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sys_clk_s1_arb_share_counter_next_value assignment, which is an e_assign
  sys_clk_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sys_clk_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sys_clk_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sys_clk_s1_allgrants all slave grants, which is an e_mux
  sys_clk_s1_allgrants <= sys_clk_s1_grant_vector;
  --sys_clk_s1_end_xfer assignment, which is an e_assign
  sys_clk_s1_end_xfer <= NOT ((sys_clk_s1_waits_for_read OR sys_clk_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sys_clk_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sys_clk_s1 <= sys_clk_s1_end_xfer AND (((NOT sys_clk_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sys_clk_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sys_clk_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sys_clk_s1 AND sys_clk_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sys_clk_s1 AND NOT sys_clk_s1_non_bursting_master_requests));
  --sys_clk_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sys_clk_s1_arb_counter_enable) = '1' then 
        sys_clk_s1_arb_share_counter <= sys_clk_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sys_clk_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sys_clk_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_sys_clk_s1)) OR ((end_xfer_arb_share_counter_term_sys_clk_s1 AND NOT sys_clk_s1_non_bursting_master_requests)))) = '1' then 
        sys_clk_s1_slavearbiterlockenable <= sys_clk_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 sys_clk/s1 arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= sys_clk_s1_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --sys_clk_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sys_clk_s1_slavearbiterlockenable2 <= sys_clk_s1_arb_share_counter_next_value;
  --clock_crossing_0/m1 sys_clk/s1 arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= sys_clk_s1_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --sys_clk_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  sys_clk_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_sys_clk_s1 <= internal_clock_crossing_0_m1_requests_sys_clk_s1 AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_sys_clk_s1, which is an e_mux
  clock_crossing_0_m1_read_data_valid_sys_clk_s1 <= (internal_clock_crossing_0_m1_granted_sys_clk_s1 AND clock_crossing_0_m1_read) AND NOT sys_clk_s1_waits_for_read;
  --sys_clk_s1_writedata mux, which is an e_mux
  sys_clk_s1_writedata <= clock_crossing_0_m1_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_sys_clk_s1 <= internal_clock_crossing_0_m1_qualified_request_sys_clk_s1;
  --clock_crossing_0/m1 saved-grant sys_clk/s1, which is an e_assign
  clock_crossing_0_m1_saved_grant_sys_clk_s1 <= internal_clock_crossing_0_m1_requests_sys_clk_s1;
  --allow new arb cycle for sys_clk/s1, which is an e_assign
  sys_clk_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sys_clk_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sys_clk_s1_master_qreq_vector <= std_logic'('1');
  --sys_clk_s1_reset_n assignment, which is an e_assign
  sys_clk_s1_reset_n <= reset_n;
  sys_clk_s1_chipselect <= internal_clock_crossing_0_m1_granted_sys_clk_s1;
  --sys_clk_s1_firsttransfer first transaction, which is an e_assign
  sys_clk_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sys_clk_s1_begins_xfer) = '1'), sys_clk_s1_unreg_firsttransfer, sys_clk_s1_reg_firsttransfer);
  --sys_clk_s1_unreg_firsttransfer first transaction, which is an e_assign
  sys_clk_s1_unreg_firsttransfer <= NOT ((sys_clk_s1_slavearbiterlockenable AND sys_clk_s1_any_continuerequest));
  --sys_clk_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sys_clk_s1_begins_xfer) = '1' then 
        sys_clk_s1_reg_firsttransfer <= sys_clk_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sys_clk_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sys_clk_s1_beginbursttransfer_internal <= sys_clk_s1_begins_xfer;
  --~sys_clk_s1_write_n assignment, which is an e_mux
  sys_clk_s1_write_n <= NOT ((internal_clock_crossing_0_m1_granted_sys_clk_s1 AND clock_crossing_0_m1_write));
  --sys_clk_s1_address mux, which is an e_mux
  sys_clk_s1_address <= clock_crossing_0_m1_nativeaddress (2 DOWNTO 0);
  --d1_sys_clk_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sys_clk_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sys_clk_s1_end_xfer <= sys_clk_s1_end_xfer;
    end if;

  end process;

  --sys_clk_s1_waits_for_read in a cycle, which is an e_mux
  sys_clk_s1_waits_for_read <= sys_clk_s1_in_a_read_cycle AND sys_clk_s1_begins_xfer;
  --sys_clk_s1_in_a_read_cycle assignment, which is an e_assign
  sys_clk_s1_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_sys_clk_s1 AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sys_clk_s1_in_a_read_cycle;
  --sys_clk_s1_waits_for_write in a cycle, which is an e_mux
  sys_clk_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sys_clk_s1_in_a_write_cycle assignment, which is an e_assign
  sys_clk_s1_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_sys_clk_s1 AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sys_clk_s1_in_a_write_cycle;
  wait_for_sys_clk_s1_counter <= std_logic'('0');
  --assign sys_clk_s1_irq_from_sa = sys_clk_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sys_clk_s1_irq_from_sa <= sys_clk_s1_irq;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_sys_clk_s1 <= internal_clock_crossing_0_m1_granted_sys_clk_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_sys_clk_s1 <= internal_clock_crossing_0_m1_qualified_request_sys_clk_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_sys_clk_s1 <= internal_clock_crossing_0_m1_requests_sys_clk_s1;
--synthesis translate_off
    --sys_clk/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_edm1_reset_cpu_clk_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity gpib_edm1_reset_cpu_clk_domain_synch_module;


architecture europa of gpib_edm1_reset_cpu_clk_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_edm1_reset_ddr_sdram_phy_clk_out_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity gpib_edm1_reset_ddr_sdram_phy_clk_out_domain_synch_module;


architecture europa of gpib_edm1_reset_ddr_sdram_phy_clk_out_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_edm1_reset_pll_c2_out_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity gpib_edm1_reset_pll_c2_out_domain_synch_module;


architecture europa of gpib_edm1_reset_pll_c2_out_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_edm1_reset_pll_c3_out_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity gpib_edm1_reset_pll_c3_out_domain_synch_module;


architecture europa of gpib_edm1_reset_pll_c3_out_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity gpib_edm1 is 
        port (
              -- 1) global signals:
                 signal clk_0 : IN STD_LOGIC;
                 signal cpu_clk : OUT STD_LOGIC;
                 signal ddr_sdram_aux_full_rate_clk_out : OUT STD_LOGIC;
                 signal ddr_sdram_aux_half_rate_clk_out : OUT STD_LOGIC;
                 signal ddr_sdram_phy_clk_out : OUT STD_LOGIC;
                 signal pll_c2_out : OUT STD_LOGIC;
                 signal pll_c3_out : OUT STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal ssram_clk : OUT STD_LOGIC;

              -- the_ad7928
                 signal MISO_to_the_ad7928 : IN STD_LOGIC;
                 signal MOSI_from_the_ad7928 : OUT STD_LOGIC;
                 signal SCLK_from_the_ad7928 : OUT STD_LOGIC;
                 signal SS_n_from_the_ad7928 : OUT STD_LOGIC;

              -- the_dac_ad5308
                 signal MISO_to_the_dac_ad5308 : IN STD_LOGIC;
                 signal MOSI_from_the_dac_ad5308 : OUT STD_LOGIC;
                 signal SCLK_from_the_dac_ad5308 : OUT STD_LOGIC;
                 signal SS_n_from_the_dac_ad5308 : OUT STD_LOGIC;

              -- the_ddr_sdram
                 signal global_reset_n_to_the_ddr_sdram : IN STD_LOGIC;
                 signal local_init_done_from_the_ddr_sdram : OUT STD_LOGIC;
                 signal local_refresh_ack_from_the_ddr_sdram : OUT STD_LOGIC;
                 signal local_wdata_req_from_the_ddr_sdram : OUT STD_LOGIC;
                 signal mem_addr_from_the_ddr_sdram : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal mem_ba_from_the_ddr_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal mem_cas_n_from_the_ddr_sdram : OUT STD_LOGIC;
                 signal mem_cke_from_the_ddr_sdram : OUT STD_LOGIC;
                 signal mem_clk_n_to_and_from_the_ddr_sdram : INOUT STD_LOGIC;
                 signal mem_clk_to_and_from_the_ddr_sdram : INOUT STD_LOGIC;
                 signal mem_cs_n_from_the_ddr_sdram : OUT STD_LOGIC;
                 signal mem_dm_from_the_ddr_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal mem_dq_to_and_from_the_ddr_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal mem_dqs_to_and_from_the_ddr_sdram : INOUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal mem_ras_n_from_the_ddr_sdram : OUT STD_LOGIC;
                 signal mem_we_n_from_the_ddr_sdram : OUT STD_LOGIC;
                 signal reset_phy_clk_n_from_the_ddr_sdram : OUT STD_LOGIC;

              -- the_flash_ssram_tristate_avalon_slave
                 signal adsc_n_to_the_ssram : OUT STD_LOGIC;
                 signal bw_n_to_the_ssram : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal bwe_n_to_the_ssram : OUT STD_LOGIC;
                 signal chipenable1_n_to_the_ssram : OUT STD_LOGIC;
                 signal flash_ssram_tristate_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal flash_ssram_tristate_data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal outputenable_n_to_the_ssram : OUT STD_LOGIC;
                 signal read_n_to_the_cfi_flash : OUT STD_LOGIC;
                 signal reset_n_to_the_ssram : OUT STD_LOGIC;
                 signal select_n_to_the_cfi_flash : OUT STD_LOGIC;
                 signal write_n_to_the_cfi_flash : OUT STD_LOGIC;

              -- the_gpib_leds
                 signal out_port_from_the_gpib_leds : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_gpio1
                 signal bidir_port_to_and_from_the_gpio1 : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_gpio2
                 signal out_port_from_the_gpio2 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_led_pio
                 signal out_port_from_the_led_pio : OUT STD_LOGIC
              );
end entity gpib_edm1;


architecture europa of gpib_edm1 is
component ad7928_spi_control_port_arbitrator is 
           port (
                 -- inputs:
                    signal ad7928_spi_control_port_dataavailable : IN STD_LOGIC;
                    signal ad7928_spi_control_port_endofpacket : IN STD_LOGIC;
                    signal ad7928_spi_control_port_irq : IN STD_LOGIC;
                    signal ad7928_spi_control_port_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal ad7928_spi_control_port_readyfordata : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_2_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal gpib_edm1_clock_2_out_read : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_out_write : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal ad7928_spi_control_port_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal ad7928_spi_control_port_chipselect : OUT STD_LOGIC;
                    signal ad7928_spi_control_port_dataavailable_from_sa : OUT STD_LOGIC;
                    signal ad7928_spi_control_port_endofpacket_from_sa : OUT STD_LOGIC;
                    signal ad7928_spi_control_port_irq_from_sa : OUT STD_LOGIC;
                    signal ad7928_spi_control_port_read_n : OUT STD_LOGIC;
                    signal ad7928_spi_control_port_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal ad7928_spi_control_port_readyfordata_from_sa : OUT STD_LOGIC;
                    signal ad7928_spi_control_port_reset_n : OUT STD_LOGIC;
                    signal ad7928_spi_control_port_write_n : OUT STD_LOGIC;
                    signal ad7928_spi_control_port_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal d1_ad7928_spi_control_port_end_xfer : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_out_granted_ad7928_spi_control_port : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_out_read_data_valid_ad7928_spi_control_port : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_out_requests_ad7928_spi_control_port : OUT STD_LOGIC
                 );
end component ad7928_spi_control_port_arbitrator;

component ad7928 is 
           port (
                 -- inputs:
                    signal MISO : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_from_cpu : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal mem_addr : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal read_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal spi_select : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;

                 -- outputs:
                    signal MOSI : OUT STD_LOGIC;
                    signal SCLK : OUT STD_LOGIC;
                    signal SS_n : OUT STD_LOGIC;
                    signal data_to_cpu : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal dataavailable : OUT STD_LOGIC;
                    signal endofpacket : OUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component ad7928;

component clock_crossing_0_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_s1_endofpacket : IN STD_LOGIC;
                    signal clock_crossing_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_0_s1_readdatavalid : IN STD_LOGIC;
                    signal clock_crossing_0_s1_waitrequest : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_instruction_master_read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_s1_address : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_0_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal clock_crossing_0_s1_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_s1_read : OUT STD_LOGIC;
                    signal clock_crossing_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_0_s1_reset_n : OUT STD_LOGIC;
                    signal clock_crossing_0_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal clock_crossing_0_s1_write : OUT STD_LOGIC;
                    signal clock_crossing_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_data_master_granted_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_granted_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_requests_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal d1_clock_crossing_0_s1_end_xfer : OUT STD_LOGIC
                 );
end component clock_crossing_0_s1_arbitrator;

component clock_crossing_0_m1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_0_m1_granted_gpib_edm1_clock_2_in : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_gpib_edm1_clock_3_in : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_gpib_leds_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_gpio1_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_gpio2_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_high_res_timer_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_led_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_sys_clk_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_gpib_leds_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_gpio1_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_gpio2_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_high_res_timer_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_led_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_sys_clk_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_gpib_leds_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_gpio1_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_gpio2_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_high_res_timer_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_led_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_sys_clk_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_gpib_edm1_clock_2_in : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_gpib_edm1_clock_3_in : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_gpib_leds_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_gpio1_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_gpio2_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_high_res_timer_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_led_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_sys_clk_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_gpib_edm1_clock_2_in_end_xfer : IN STD_LOGIC;
                    signal d1_gpib_edm1_clock_3_in_end_xfer : IN STD_LOGIC;
                    signal d1_gpib_leds_s1_end_xfer : IN STD_LOGIC;
                    signal d1_gpio1_s1_end_xfer : IN STD_LOGIC;
                    signal d1_gpio2_s1_end_xfer : IN STD_LOGIC;
                    signal d1_high_res_timer_s1_end_xfer : IN STD_LOGIC;
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                    signal d1_led_pio_s1_end_xfer : IN STD_LOGIC;
                    signal d1_sys_clk_s1_end_xfer : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_in_endofpacket_from_sa : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_2_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_in_endofpacket_from_sa : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_3_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal gpib_leds_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gpio1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gpio2_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal high_res_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal led_pio_s1_readdata_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal clock_crossing_0_m1_address_to_slave : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_endofpacket : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_latency_counter : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_0_m1_readdatavalid : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_reset_n : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_waitrequest : OUT STD_LOGIC
                 );
end component clock_crossing_0_m1_arbitrator;

component clock_crossing_0 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_readdatavalid : IN STD_LOGIC;
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_readdatavalid : OUT STD_LOGIC;
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component clock_crossing_0;

component clock_crossing_0_bridge_arbitrator is 
end component clock_crossing_0_bridge_arbitrator;

component cpu_0_jtag_debug_module_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_instruction_master_read : IN STD_LOGIC;
                    signal cpu_0_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_jtag_debug_module_resetrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_granted_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_requests_cpu_0_jtag_debug_module : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal cpu_0_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_jtag_debug_module_chipselect : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_jtag_debug_module_reset_n : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_write : OUT STD_LOGIC;
                    signal cpu_0_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_0_jtag_debug_module_end_xfer : OUT STD_LOGIC
                 );
end component cpu_0_jtag_debug_module_arbitrator;

component cpu_0_data_master_arbitrator is 
           port (
                 -- inputs:
                    signal ad7928_spi_control_port_irq_from_sa : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_0_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal cpu_0_data_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_data_master_granted_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_gpib_edm1_clock_0_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_gpib_edm1_clock_1_in : IN STD_LOGIC;
                    signal cpu_0_data_master_granted_onchip_memory_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in : IN STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_onchip_memory_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_gpib_edm1_clock_0_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_gpib_edm1_clock_1_in : IN STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_onchip_memory_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_gpib_edm1_clock_0_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_gpib_edm1_clock_1_in : IN STD_LOGIC;
                    signal cpu_0_data_master_requests_onchip_memory_s1 : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_clk : IN STD_LOGIC;
                    signal cpu_clk_reset_n : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal d1_clock_crossing_0_s1_end_xfer : IN STD_LOGIC;
                    signal d1_cpu_0_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_cpu_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal d1_flash_ssram_pipeline_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal d1_gpib_edm1_clock_0_in_end_xfer : IN STD_LOGIC;
                    signal d1_gpib_edm1_clock_1_in_end_xfer : IN STD_LOGIC;
                    signal d1_onchip_memory_s1_end_xfer : IN STD_LOGIC;
                    signal dac_ad5308_spi_control_port_irq_from_sa : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpib_edm1_clock_1_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal high_res_timer_s1_irq_from_sa : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                    signal onchip_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal registered_cpu_0_data_master_read_data_valid_onchip_memory_s1 : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_s1_irq_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_data_master_waitrequest : OUT STD_LOGIC
                 );
end component cpu_0_data_master_arbitrator;

component cpu_0_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_0_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal cpu_0_instruction_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_instruction_master_granted_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_granted_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_granted_onchip_memory_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_onchip_memory_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_onchip_memory_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_requests_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_requests_cpu_0_jtag_debug_module : IN STD_LOGIC;
                    signal cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_0_instruction_master_requests_onchip_memory_s1 : IN STD_LOGIC;
                    signal cpu_0_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal d1_clock_crossing_0_s1_end_xfer : IN STD_LOGIC;
                    signal d1_cpu_0_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_cpu_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal d1_flash_ssram_pipeline_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal d1_onchip_memory_s1_end_xfer : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal onchip_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_instruction_master_waitrequest : OUT STD_LOGIC
                 );
end component cpu_0_instruction_master_arbitrator;

component cpu_0 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d_irq : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_waitrequest : IN STD_LOGIC;
                    signal i_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_waitrequest : IN STD_LOGIC;
                    signal jtag_debug_module_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal jtag_debug_module_begintransfer : IN STD_LOGIC;
                    signal jtag_debug_module_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal jtag_debug_module_debugaccess : IN STD_LOGIC;
                    signal jtag_debug_module_select : IN STD_LOGIC;
                    signal jtag_debug_module_write : IN STD_LOGIC;
                    signal jtag_debug_module_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d_address : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal d_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_read : OUT STD_LOGIC;
                    signal d_write : OUT STD_LOGIC;
                    signal d_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_address : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal i_read : OUT STD_LOGIC;
                    signal jtag_debug_module_debugaccess_to_roms : OUT STD_LOGIC;
                    signal jtag_debug_module_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_debug_module_resetrequest : OUT STD_LOGIC
                 );
end component cpu_0;

component cpu_ddr_clock_bridge_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_instruction_master_read : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_endofpacket : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_readdatavalid : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_read : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_reset_n : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_write : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_ddr_clock_bridge_s1_end_xfer : OUT STD_LOGIC
                 );
end component cpu_ddr_clock_bridge_s1_arbitrator;

component cpu_ddr_clock_bridge_m1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1 : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1_shift_register : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_ddr_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal ddr_sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ddr_sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_ddr_clock_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_latency_counter : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_readdatavalid : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_reset_n : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_waitrequest : OUT STD_LOGIC
                 );
end component cpu_ddr_clock_bridge_m1_arbitrator;

component cpu_ddr_clock_bridge is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_readdatavalid : IN STD_LOGIC;
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_readdatavalid : OUT STD_LOGIC;
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component cpu_ddr_clock_bridge;

component cpu_ddr_clock_bridge_bridge_arbitrator is 
end component cpu_ddr_clock_bridge_bridge_arbitrator;

component dac_ad5308_spi_control_port_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal dac_ad5308_spi_control_port_dataavailable : IN STD_LOGIC;
                    signal dac_ad5308_spi_control_port_endofpacket : IN STD_LOGIC;
                    signal dac_ad5308_spi_control_port_irq : IN STD_LOGIC;
                    signal dac_ad5308_spi_control_port_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal dac_ad5308_spi_control_port_readyfordata : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_3_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal gpib_edm1_clock_3_out_read : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_out_write : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_dac_ad5308_spi_control_port_end_xfer : OUT STD_LOGIC;
                    signal dac_ad5308_spi_control_port_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal dac_ad5308_spi_control_port_chipselect : OUT STD_LOGIC;
                    signal dac_ad5308_spi_control_port_dataavailable_from_sa : OUT STD_LOGIC;
                    signal dac_ad5308_spi_control_port_endofpacket_from_sa : OUT STD_LOGIC;
                    signal dac_ad5308_spi_control_port_irq_from_sa : OUT STD_LOGIC;
                    signal dac_ad5308_spi_control_port_read_n : OUT STD_LOGIC;
                    signal dac_ad5308_spi_control_port_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal dac_ad5308_spi_control_port_readyfordata_from_sa : OUT STD_LOGIC;
                    signal dac_ad5308_spi_control_port_reset_n : OUT STD_LOGIC;
                    signal dac_ad5308_spi_control_port_write_n : OUT STD_LOGIC;
                    signal dac_ad5308_spi_control_port_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_out_read_data_valid_dac_ad5308_spi_control_port : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port : OUT STD_LOGIC
                 );
end component dac_ad5308_spi_control_port_arbitrator;

component dac_ad5308 is 
           port (
                 -- inputs:
                    signal MISO : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_from_cpu : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal mem_addr : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal read_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal spi_select : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;

                 -- outputs:
                    signal MOSI : OUT STD_LOGIC;
                    signal SCLK : OUT STD_LOGIC;
                    signal SS_n : OUT STD_LOGIC;
                    signal data_to_cpu : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal dataavailable : OUT STD_LOGIC;
                    signal endofpacket : OUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component dac_ad5308;

component ddr_sdram_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ddr_sdram_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ddr_sdram_s1_readdatavalid : IN STD_LOGIC;
                    signal ddr_sdram_s1_resetrequest_n : IN STD_LOGIC;
                    signal ddr_sdram_s1_waitrequest_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1 : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 : OUT STD_LOGIC;
                    signal d1_ddr_sdram_s1_end_xfer : OUT STD_LOGIC;
                    signal ddr_sdram_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal ddr_sdram_s1_beginbursttransfer : OUT STD_LOGIC;
                    signal ddr_sdram_s1_burstcount : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal ddr_sdram_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ddr_sdram_s1_read : OUT STD_LOGIC;
                    signal ddr_sdram_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ddr_sdram_s1_resetrequest_n_from_sa : OUT STD_LOGIC;
                    signal ddr_sdram_s1_waitrequest_n_from_sa : OUT STD_LOGIC;
                    signal ddr_sdram_s1_write : OUT STD_LOGIC;
                    signal ddr_sdram_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component ddr_sdram_s1_arbitrator;

component gpib_edm1_reset_clk_0_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component gpib_edm1_reset_clk_0_domain_synch_module;

component ddr_sdram is 
           port (
                 -- inputs:
                    signal global_reset_n : IN STD_LOGIC;
                    signal local_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal local_be : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal local_burstbegin : IN STD_LOGIC;
                    signal local_read_req : IN STD_LOGIC;
                    signal local_size : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal local_wdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal local_write_req : IN STD_LOGIC;
                    signal pll_ref_clk : IN STD_LOGIC;
                    signal soft_reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal aux_full_rate_clk : OUT STD_LOGIC;
                    signal aux_half_rate_clk : OUT STD_LOGIC;
                    signal local_init_done : OUT STD_LOGIC;
                    signal local_rdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal local_rdata_valid : OUT STD_LOGIC;
                    signal local_ready : OUT STD_LOGIC;
                    signal local_refresh_ack : OUT STD_LOGIC;
                    signal local_wdata_req : OUT STD_LOGIC;
                    signal mem_addr : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal mem_ba : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_cas_n : OUT STD_LOGIC;
                    signal mem_cke : OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
                    signal mem_clk : INOUT STD_LOGIC_VECTOR (0 DOWNTO 0);
                    signal mem_clk_n : INOUT STD_LOGIC_VECTOR (0 DOWNTO 0);
                    signal mem_cs_n : OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
                    signal mem_dm : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_dq : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal mem_dqs : INOUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_ras_n : OUT STD_LOGIC;
                    signal mem_we_n : OUT STD_LOGIC;
                    signal phy_clk : OUT STD_LOGIC;
                    signal reset_phy_clk_n : OUT STD_LOGIC;
                    signal reset_request_n : OUT STD_LOGIC
                 );
end component ddr_sdram;

component flash_ssram_pipeline_bridge_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_instruction_master_read : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_endofpacket : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_s1_readdatavalid : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal d1_flash_ssram_pipeline_bridge_s1_end_xfer : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_s1_arbiterlock : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_arbiterlock2 : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_burstcount : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_s1_chipselect : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_debugaccess : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_s1_read : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_s1_reset_n : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_write : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component flash_ssram_pipeline_bridge_s1_arbitrator;

component flash_ssram_pipeline_bridge_m1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_pipeline_bridge_before_tristate_s1_end_xfer : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1 : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1_shift_register : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_s1_endofpacket_from_sa : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal flash_ssram_pipeline_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_m1_endofpacket : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_latency_counter : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_m1_readdatavalid : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_waitrequest : OUT STD_LOGIC
                 );
end component flash_ssram_pipeline_bridge_m1_arbitrator;

component flash_ssram_pipeline_bridge is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal m1_endofpacket : IN STD_LOGIC;
                    signal m1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m1_readdatavalid : IN STD_LOGIC;
                    signal m1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal s1_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal s1_arbiterlock : IN STD_LOGIC;
                    signal s1_arbiterlock2 : IN STD_LOGIC;
                    signal s1_burstcount : IN STD_LOGIC;
                    signal s1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal s1_chipselect : IN STD_LOGIC;
                    signal s1_debugaccess : IN STD_LOGIC;
                    signal s1_nativeaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal s1_read : IN STD_LOGIC;
                    signal s1_write : IN STD_LOGIC;
                    signal s1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal m1_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal m1_burstcount : OUT STD_LOGIC;
                    signal m1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m1_chipselect : OUT STD_LOGIC;
                    signal m1_debugaccess : OUT STD_LOGIC;
                    signal m1_read : OUT STD_LOGIC;
                    signal m1_write : OUT STD_LOGIC;
                    signal m1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal s1_endofpacket : OUT STD_LOGIC;
                    signal s1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal s1_readdatavalid : OUT STD_LOGIC;
                    signal s1_waitrequest : OUT STD_LOGIC
                 );
end component flash_ssram_pipeline_bridge;

component flash_ssram_pipeline_bridge_bridge_arbitrator is 
end component flash_ssram_pipeline_bridge_bridge_arbitrator;

component flash_ssram_tristate_avalon_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal adsc_n_to_the_ssram : OUT STD_LOGIC;
                    signal bw_n_to_the_ssram : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal bwe_n_to_the_ssram : OUT STD_LOGIC;
                    signal cfi_flash_s1_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal chipenable1_n_to_the_ssram : OUT STD_LOGIC;
                    signal d1_flash_ssram_tristate_avalon_slave_end_xfer : OUT STD_LOGIC;
                    signal flash_ssram_tristate_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal flash_ssram_tristate_data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal incoming_flash_ssram_tristate_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal incoming_flash_ssram_tristate_data_with_Xs_converted_to_0 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal outputenable_n_to_the_ssram : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_granted_ssram_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_requests_ssram_s1 : OUT STD_LOGIC;
                    signal read_n_to_the_cfi_flash : OUT STD_LOGIC;
                    signal reset_n_to_the_ssram : OUT STD_LOGIC;
                    signal select_n_to_the_cfi_flash : OUT STD_LOGIC;
                    signal write_n_to_the_cfi_flash : OUT STD_LOGIC
                 );
end component flash_ssram_tristate_avalon_slave_arbitrator;

component flash_ssram_tristate is 
end component flash_ssram_tristate;

component flash_ssram_tristate_bridge_arbitrator is 
end component flash_ssram_tristate_bridge_arbitrator;

component gpib_edm1_clock_0_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpib_edm1_clock_0_in_endofpacket : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_0_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_gpib_edm1_clock_0_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_gpib_edm1_clock_0_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_gpib_edm1_clock_0_in : OUT STD_LOGIC;
                    signal d1_gpib_edm1_clock_0_in_end_xfer : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gpib_edm1_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal gpib_edm1_clock_0_in_read : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_0_in_reset_n : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_in_write : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component gpib_edm1_clock_0_in_arbitrator;

component gpib_edm1_clock_0_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_pll_s1_end_xfer : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gpib_edm1_clock_0_out_granted_pll_s1 : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_out_qualified_request_pll_s1 : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_out_read : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_out_read_data_valid_pll_s1 : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_out_requests_pll_s1 : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_out_write : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pll_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal gpib_edm1_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_0_out_reset_n : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_out_waitrequest : OUT STD_LOGIC
                 );
end component gpib_edm1_clock_0_out_arbitrator;

component gpib_edm1_clock_0 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component gpib_edm1_clock_0;

component gpib_edm1_clock_1_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpib_edm1_clock_1_in_endofpacket : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpib_edm1_clock_1_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_gpib_edm1_clock_1_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_gpib_edm1_clock_1_in : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_gpib_edm1_clock_1_in : OUT STD_LOGIC;
                    signal d1_gpib_edm1_clock_1_in_end_xfer : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_in_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gpib_edm1_clock_1_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_1_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_in_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal gpib_edm1_clock_1_in_read : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpib_edm1_clock_1_in_reset_n : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_in_write : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component gpib_edm1_clock_1_in_arbitrator;

component gpib_edm1_clock_1_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_remote_update_cycloneiii_1_s1_end_xfer : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_out_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gpib_edm1_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_out_read : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1 : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_out_write : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal remote_update_cycloneiii_1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal remote_update_cycloneiii_1_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal gpib_edm1_clock_1_out_address_to_slave : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gpib_edm1_clock_1_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpib_edm1_clock_1_out_reset_n : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_out_waitrequest : OUT STD_LOGIC
                 );
end component gpib_edm1_clock_1_out_arbitrator;

component gpib_edm1_clock_1 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component gpib_edm1_clock_1;

component gpib_edm1_clock_2_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpib_edm1_clock_2_in_endofpacket : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_2_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_m1_granted_gpib_edm1_clock_2_in : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_gpib_edm1_clock_2_in : OUT STD_LOGIC;
                    signal d1_gpib_edm1_clock_2_in_end_xfer : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_2_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gpib_edm1_clock_2_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal gpib_edm1_clock_2_in_read : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_2_in_reset_n : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_in_write : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component gpib_edm1_clock_2_in_arbitrator;

component gpib_edm1_clock_2_out_arbitrator is 
           port (
                 -- inputs:
                    signal ad7928_spi_control_port_endofpacket_from_sa : IN STD_LOGIC;
                    signal ad7928_spi_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_ad7928_spi_control_port_end_xfer : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_2_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gpib_edm1_clock_2_out_granted_ad7928_spi_control_port : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_out_read : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_out_read_data_valid_ad7928_spi_control_port : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_out_requests_ad7928_spi_control_port : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_out_write : IN STD_LOGIC;
                    signal gpib_edm1_clock_2_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal gpib_edm1_clock_2_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_2_out_endofpacket : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_2_out_reset_n : OUT STD_LOGIC;
                    signal gpib_edm1_clock_2_out_waitrequest : OUT STD_LOGIC
                 );
end component gpib_edm1_clock_2_out_arbitrator;

component gpib_edm1_clock_2 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component gpib_edm1_clock_2;

component gpib_edm1_clock_3_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpib_edm1_clock_3_in_endofpacket : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_3_in_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_m1_granted_gpib_edm1_clock_3_in : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_gpib_edm1_clock_3_in : OUT STD_LOGIC;
                    signal d1_gpib_edm1_clock_3_in_end_xfer : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_3_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gpib_edm1_clock_3_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal gpib_edm1_clock_3_in_read : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_3_in_reset_n : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_in_write : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component gpib_edm1_clock_3_in_arbitrator;

component gpib_edm1_clock_3_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_dac_ad5308_spi_control_port_end_xfer : IN STD_LOGIC;
                    signal dac_ad5308_spi_control_port_endofpacket_from_sa : IN STD_LOGIC;
                    signal dac_ad5308_spi_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_3_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_3_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_out_read : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_out_read_data_valid_dac_ad5308_spi_control_port : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_out_write : IN STD_LOGIC;
                    signal gpib_edm1_clock_3_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal gpib_edm1_clock_3_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_3_out_endofpacket : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal gpib_edm1_clock_3_out_reset_n : OUT STD_LOGIC;
                    signal gpib_edm1_clock_3_out_waitrequest : OUT STD_LOGIC
                 );
end component gpib_edm1_clock_3_out_arbitrator;

component gpib_edm1_clock_3 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component gpib_edm1_clock_3;

component gpib_leds_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpib_leds_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_m1_granted_gpib_leds_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_gpib_leds_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_gpib_leds_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_gpib_leds_s1 : OUT STD_LOGIC;
                    signal d1_gpib_leds_s1_end_xfer : OUT STD_LOGIC;
                    signal gpib_leds_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gpib_leds_s1_chipselect : OUT STD_LOGIC;
                    signal gpib_leds_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gpib_leds_s1_reset_n : OUT STD_LOGIC;
                    signal gpib_leds_s1_write_n : OUT STD_LOGIC;
                    signal gpib_leds_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component gpib_leds_s1_arbitrator;

component gpib_leds is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component gpib_leds;

component gpio1_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpio1_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_m1_granted_gpio1_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_gpio1_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_gpio1_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_gpio1_s1 : OUT STD_LOGIC;
                    signal d1_gpio1_s1_end_xfer : OUT STD_LOGIC;
                    signal gpio1_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal gpio1_s1_chipselect : OUT STD_LOGIC;
                    signal gpio1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gpio1_s1_reset_n : OUT STD_LOGIC;
                    signal gpio1_s1_write_n : OUT STD_LOGIC;
                    signal gpio1_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component gpio1_s1_arbitrator;

component gpio1 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal bidir_port : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component gpio1;

component gpio2_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal gpio2_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_m1_granted_gpio2_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_gpio2_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_gpio2_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_gpio2_s1 : OUT STD_LOGIC;
                    signal d1_gpio2_s1_end_xfer : OUT STD_LOGIC;
                    signal gpio2_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal gpio2_s1_chipselect : OUT STD_LOGIC;
                    signal gpio2_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gpio2_s1_reset_n : OUT STD_LOGIC;
                    signal gpio2_s1_write_n : OUT STD_LOGIC;
                    signal gpio2_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component gpio2_s1_arbitrator;

component gpio2 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component gpio2;

component high_res_timer_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal high_res_timer_s1_irq : IN STD_LOGIC;
                    signal high_res_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_m1_granted_high_res_timer_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_high_res_timer_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_high_res_timer_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_high_res_timer_s1 : OUT STD_LOGIC;
                    signal d1_high_res_timer_s1_end_xfer : OUT STD_LOGIC;
                    signal high_res_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal high_res_timer_s1_chipselect : OUT STD_LOGIC;
                    signal high_res_timer_s1_irq_from_sa : OUT STD_LOGIC;
                    signal high_res_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal high_res_timer_s1_reset_n : OUT STD_LOGIC;
                    signal high_res_timer_s1_write_n : OUT STD_LOGIC;
                    signal high_res_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component high_res_timer_s1_arbitrator;

component high_res_timer is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component high_res_timer;

component jtag_uart_avalon_jtag_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component jtag_uart_avalon_jtag_slave_arbitrator;

component jtag_uart is 
           port (
                 -- inputs:
                    signal av_address : IN STD_LOGIC;
                    signal av_chipselect : IN STD_LOGIC;
                    signal av_read_n : IN STD_LOGIC;
                    signal av_write_n : IN STD_LOGIC;
                    signal av_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_irq : OUT STD_LOGIC;
                    signal av_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_waitrequest : OUT STD_LOGIC;
                    signal dataavailable : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component jtag_uart;

component led_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal led_pio_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_m1_granted_led_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_led_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_led_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_led_pio_s1 : OUT STD_LOGIC;
                    signal d1_led_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal led_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal led_pio_s1_chipselect : OUT STD_LOGIC;
                    signal led_pio_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal led_pio_s1_reset_n : OUT STD_LOGIC;
                    signal led_pio_s1_write_n : OUT STD_LOGIC;
                    signal led_pio_s1_writedata : OUT STD_LOGIC
                 );
end component led_pio_s1_arbitrator;

component led_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component led_pio;

component onchip_memory_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_0_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_0_data_master_read : IN STD_LOGIC;
                    signal cpu_0_data_master_waitrequest : IN STD_LOGIC;
                    signal cpu_0_data_master_write : IN STD_LOGIC;
                    signal cpu_0_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_0_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_0_instruction_master_read : IN STD_LOGIC;
                    signal onchip_memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_0_data_master_granted_onchip_memory_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_qualified_request_onchip_memory_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_read_data_valid_onchip_memory_s1 : OUT STD_LOGIC;
                    signal cpu_0_data_master_requests_onchip_memory_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_granted_onchip_memory_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_qualified_request_onchip_memory_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_read_data_valid_onchip_memory_s1 : OUT STD_LOGIC;
                    signal cpu_0_instruction_master_requests_onchip_memory_s1 : OUT STD_LOGIC;
                    signal d1_onchip_memory_s1_end_xfer : OUT STD_LOGIC;
                    signal onchip_memory_s1_address : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal onchip_memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal onchip_memory_s1_chipselect : OUT STD_LOGIC;
                    signal onchip_memory_s1_clken : OUT STD_LOGIC;
                    signal onchip_memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal onchip_memory_s1_reset : OUT STD_LOGIC;
                    signal onchip_memory_s1_write : OUT STD_LOGIC;
                    signal onchip_memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal registered_cpu_0_data_master_read_data_valid_onchip_memory_s1 : OUT STD_LOGIC
                 );
end component onchip_memory_s1_arbitrator;

component onchip_memory is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clken : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component onchip_memory;

component pipeline_bridge_before_tristate_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal flash_ssram_pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_debugaccess : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_s1_endofpacket : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_s1_readdatavalid : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pipeline_bridge_before_tristate_s1_end_xfer : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1 : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1_shift_register : OUT STD_LOGIC;
                    signal flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_s1_arbiterlock : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_arbiterlock2 : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_burstcount : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_s1_chipselect : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_debugaccess : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_s1_read : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_s1_reset_n : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_write : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component pipeline_bridge_before_tristate_s1_arbitrator;

component pipeline_bridge_before_tristate_m1_arbitrator is 
           port (
                 -- inputs:
                    signal cfi_flash_s1_wait_counter_eq_0 : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal d1_flash_ssram_tristate_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal incoming_flash_ssram_tristate_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal incoming_flash_ssram_tristate_data_with_Xs_converted_to_0 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_granted_ssram_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_requests_ssram_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal pipeline_bridge_before_tristate_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_latency_counter : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_before_tristate_m1_readdatavalid : OUT STD_LOGIC;
                    signal pipeline_bridge_before_tristate_m1_waitrequest : OUT STD_LOGIC
                 );
end component pipeline_bridge_before_tristate_m1_arbitrator;

component pipeline_bridge_before_tristate is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal m1_endofpacket : IN STD_LOGIC;
                    signal m1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m1_readdatavalid : IN STD_LOGIC;
                    signal m1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal s1_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal s1_arbiterlock : IN STD_LOGIC;
                    signal s1_arbiterlock2 : IN STD_LOGIC;
                    signal s1_burstcount : IN STD_LOGIC;
                    signal s1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal s1_chipselect : IN STD_LOGIC;
                    signal s1_debugaccess : IN STD_LOGIC;
                    signal s1_nativeaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal s1_read : IN STD_LOGIC;
                    signal s1_write : IN STD_LOGIC;
                    signal s1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal m1_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal m1_burstcount : OUT STD_LOGIC;
                    signal m1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m1_chipselect : OUT STD_LOGIC;
                    signal m1_debugaccess : OUT STD_LOGIC;
                    signal m1_read : OUT STD_LOGIC;
                    signal m1_write : OUT STD_LOGIC;
                    signal m1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal s1_endofpacket : OUT STD_LOGIC;
                    signal s1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal s1_readdatavalid : OUT STD_LOGIC;
                    signal s1_waitrequest : OUT STD_LOGIC
                 );
end component pipeline_bridge_before_tristate;

component pipeline_bridge_before_tristate_bridge_arbitrator is 
end component pipeline_bridge_before_tristate_bridge_arbitrator;

component pll_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal gpib_edm1_clock_0_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal gpib_edm1_clock_0_out_read : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_out_write : IN STD_LOGIC;
                    signal gpib_edm1_clock_0_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pll_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pll_s1_resetrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pll_s1_end_xfer : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_out_granted_pll_s1 : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_out_qualified_request_pll_s1 : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_out_read_data_valid_pll_s1 : OUT STD_LOGIC;
                    signal gpib_edm1_clock_0_out_requests_pll_s1 : OUT STD_LOGIC;
                    signal pll_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal pll_s1_chipselect : OUT STD_LOGIC;
                    signal pll_s1_read : OUT STD_LOGIC;
                    signal pll_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pll_s1_reset_n : OUT STD_LOGIC;
                    signal pll_s1_resetrequest_from_sa : OUT STD_LOGIC;
                    signal pll_s1_write : OUT STD_LOGIC;
                    signal pll_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pll_s1_arbitrator;

component pll is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal c0 : OUT STD_LOGIC;
                    signal c1 : OUT STD_LOGIC;
                    signal c2 : OUT STD_LOGIC;
                    signal c3 : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal resetrequest : OUT STD_LOGIC
                 );
end component pll;

component remote_update_cycloneiii_1_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_out_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gpib_edm1_clock_1_out_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal gpib_edm1_clock_1_out_read : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_out_write : IN STD_LOGIC;
                    signal gpib_edm1_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal remote_update_cycloneiii_1_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal remote_update_cycloneiii_1_s1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_remote_update_cycloneiii_1_s1_end_xfer : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1 : OUT STD_LOGIC;
                    signal gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_1_s1_address : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal remote_update_cycloneiii_1_s1_chipselect : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_1_s1_read : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal remote_update_cycloneiii_1_s1_reset : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_1_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_1_s1_write : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_1_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component remote_update_cycloneiii_1_s1_arbitrator;

component remote_update_cycloneiii_1 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal waitrequest : OUT STD_LOGIC
                 );
end component remote_update_cycloneiii_1;

component sys_clk_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_s1_irq : IN STD_LOGIC;
                    signal sys_clk_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal clock_crossing_0_m1_granted_sys_clk_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_sys_clk_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_sys_clk_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_sys_clk_s1 : OUT STD_LOGIC;
                    signal d1_sys_clk_s1_end_xfer : OUT STD_LOGIC;
                    signal sys_clk_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal sys_clk_s1_chipselect : OUT STD_LOGIC;
                    signal sys_clk_s1_irq_from_sa : OUT STD_LOGIC;
                    signal sys_clk_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sys_clk_s1_reset_n : OUT STD_LOGIC;
                    signal sys_clk_s1_write_n : OUT STD_LOGIC;
                    signal sys_clk_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sys_clk_s1_arbitrator;

component sys_clk is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sys_clk;

component gpib_edm1_reset_cpu_clk_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component gpib_edm1_reset_cpu_clk_domain_synch_module;

component gpib_edm1_reset_ddr_sdram_phy_clk_out_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component gpib_edm1_reset_ddr_sdram_phy_clk_out_domain_synch_module;

component gpib_edm1_reset_pll_c2_out_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component gpib_edm1_reset_pll_c2_out_domain_synch_module;

component gpib_edm1_reset_pll_c3_out_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component gpib_edm1_reset_pll_c3_out_domain_synch_module;

                signal ad7928_spi_control_port_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal ad7928_spi_control_port_chipselect :  STD_LOGIC;
                signal ad7928_spi_control_port_dataavailable :  STD_LOGIC;
                signal ad7928_spi_control_port_dataavailable_from_sa :  STD_LOGIC;
                signal ad7928_spi_control_port_endofpacket :  STD_LOGIC;
                signal ad7928_spi_control_port_endofpacket_from_sa :  STD_LOGIC;
                signal ad7928_spi_control_port_irq :  STD_LOGIC;
                signal ad7928_spi_control_port_irq_from_sa :  STD_LOGIC;
                signal ad7928_spi_control_port_read_n :  STD_LOGIC;
                signal ad7928_spi_control_port_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal ad7928_spi_control_port_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal ad7928_spi_control_port_readyfordata :  STD_LOGIC;
                signal ad7928_spi_control_port_readyfordata_from_sa :  STD_LOGIC;
                signal ad7928_spi_control_port_reset_n :  STD_LOGIC;
                signal ad7928_spi_control_port_write_n :  STD_LOGIC;
                signal ad7928_spi_control_port_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal cfi_flash_s1_wait_counter_eq_0 :  STD_LOGIC;
                signal clk_0_reset_n :  STD_LOGIC;
                signal clock_crossing_0_m1_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal clock_crossing_0_m1_address_to_slave :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal clock_crossing_0_m1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clock_crossing_0_m1_endofpacket :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_gpib_edm1_clock_2_in :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_gpib_edm1_clock_3_in :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_gpib_leds_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_gpio1_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_gpio2_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_high_res_timer_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_led_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_sys_clk_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_latency_counter :  STD_LOGIC;
                signal clock_crossing_0_m1_nativeaddress :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_gpib_leds_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_gpio1_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_gpio2_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_high_res_timer_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_led_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_sys_clk_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_read :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_gpib_leds_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_gpio1_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_gpio2_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_high_res_timer_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_led_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_sys_clk_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_0_m1_readdatavalid :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_gpib_edm1_clock_2_in :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_gpib_edm1_clock_3_in :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_gpib_leds_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_gpio1_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_gpio2_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_high_res_timer_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_led_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_sys_clk_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_reset_n :  STD_LOGIC;
                signal clock_crossing_0_m1_waitrequest :  STD_LOGIC;
                signal clock_crossing_0_m1_write :  STD_LOGIC;
                signal clock_crossing_0_m1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_0_s1_address :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal clock_crossing_0_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clock_crossing_0_s1_endofpacket :  STD_LOGIC;
                signal clock_crossing_0_s1_endofpacket_from_sa :  STD_LOGIC;
                signal clock_crossing_0_s1_nativeaddress :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal clock_crossing_0_s1_read :  STD_LOGIC;
                signal clock_crossing_0_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_0_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_0_s1_readdatavalid :  STD_LOGIC;
                signal clock_crossing_0_s1_reset_n :  STD_LOGIC;
                signal clock_crossing_0_s1_waitrequest :  STD_LOGIC;
                signal clock_crossing_0_s1_waitrequest_from_sa :  STD_LOGIC;
                signal clock_crossing_0_s1_write :  STD_LOGIC;
                signal clock_crossing_0_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_data_master_address :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_0_data_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_0_data_master_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_0_data_master_debugaccess :  STD_LOGIC;
                signal cpu_0_data_master_granted_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_data_master_granted_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_granted_gpib_edm1_clock_0_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_gpib_edm1_clock_1_in :  STD_LOGIC;
                signal cpu_0_data_master_granted_onchip_memory_s1 :  STD_LOGIC;
                signal cpu_0_data_master_irq :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_data_master_qualified_request_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in :  STD_LOGIC;
                signal cpu_0_data_master_qualified_request_onchip_memory_s1 :  STD_LOGIC;
                signal cpu_0_data_master_read :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_gpib_edm1_clock_0_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_gpib_edm1_clock_1_in :  STD_LOGIC;
                signal cpu_0_data_master_read_data_valid_onchip_memory_s1 :  STD_LOGIC;
                signal cpu_0_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_data_master_requests_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_data_master_requests_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_data_master_requests_gpib_edm1_clock_0_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_gpib_edm1_clock_1_in :  STD_LOGIC;
                signal cpu_0_data_master_requests_onchip_memory_s1 :  STD_LOGIC;
                signal cpu_0_data_master_waitrequest :  STD_LOGIC;
                signal cpu_0_data_master_write :  STD_LOGIC;
                signal cpu_0_data_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_instruction_master_address :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_0_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_0_instruction_master_granted_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_granted_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_granted_onchip_memory_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_qualified_request_onchip_memory_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_read :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register :  STD_LOGIC;
                signal cpu_0_instruction_master_read_data_valid_onchip_memory_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_instruction_master_requests_clock_crossing_0_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_requests_cpu_0_jtag_debug_module :  STD_LOGIC;
                signal cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_requests_onchip_memory_s1 :  STD_LOGIC;
                signal cpu_0_instruction_master_waitrequest :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal cpu_0_jtag_debug_module_begintransfer :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_0_jtag_debug_module_chipselect :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_debugaccess :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_jtag_debug_module_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_0_jtag_debug_module_reset_n :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_resetrequest :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_resetrequest_from_sa :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_write :  STD_LOGIC;
                signal cpu_0_jtag_debug_module_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_clk_reset_n :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_endofpacket :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_latency_counter :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_read :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1_shift_register :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_readdatavalid :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_reset_n :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_waitrequest :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_write :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_endofpacket :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_read :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_readdatavalid :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_reset_n :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_waitrequest :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_write :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal d1_ad7928_spi_control_port_end_xfer :  STD_LOGIC;
                signal d1_clock_crossing_0_s1_end_xfer :  STD_LOGIC;
                signal d1_cpu_0_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal d1_cpu_ddr_clock_bridge_s1_end_xfer :  STD_LOGIC;
                signal d1_dac_ad5308_spi_control_port_end_xfer :  STD_LOGIC;
                signal d1_ddr_sdram_s1_end_xfer :  STD_LOGIC;
                signal d1_flash_ssram_pipeline_bridge_s1_end_xfer :  STD_LOGIC;
                signal d1_flash_ssram_tristate_avalon_slave_end_xfer :  STD_LOGIC;
                signal d1_gpib_edm1_clock_0_in_end_xfer :  STD_LOGIC;
                signal d1_gpib_edm1_clock_1_in_end_xfer :  STD_LOGIC;
                signal d1_gpib_edm1_clock_2_in_end_xfer :  STD_LOGIC;
                signal d1_gpib_edm1_clock_3_in_end_xfer :  STD_LOGIC;
                signal d1_gpib_leds_s1_end_xfer :  STD_LOGIC;
                signal d1_gpio1_s1_end_xfer :  STD_LOGIC;
                signal d1_gpio2_s1_end_xfer :  STD_LOGIC;
                signal d1_high_res_timer_s1_end_xfer :  STD_LOGIC;
                signal d1_jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal d1_led_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_onchip_memory_s1_end_xfer :  STD_LOGIC;
                signal d1_pipeline_bridge_before_tristate_s1_end_xfer :  STD_LOGIC;
                signal d1_pll_s1_end_xfer :  STD_LOGIC;
                signal d1_remote_update_cycloneiii_1_s1_end_xfer :  STD_LOGIC;
                signal d1_sys_clk_s1_end_xfer :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal dac_ad5308_spi_control_port_chipselect :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_dataavailable :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_dataavailable_from_sa :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_endofpacket :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_endofpacket_from_sa :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_irq :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_irq_from_sa :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_read_n :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dac_ad5308_spi_control_port_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dac_ad5308_spi_control_port_readyfordata :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_readyfordata_from_sa :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_reset_n :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_write_n :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal ddr_sdram_phy_clk_out_reset_n :  STD_LOGIC;
                signal ddr_sdram_s1_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal ddr_sdram_s1_beginbursttransfer :  STD_LOGIC;
                signal ddr_sdram_s1_burstcount :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal ddr_sdram_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_s1_read :  STD_LOGIC;
                signal ddr_sdram_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ddr_sdram_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ddr_sdram_s1_readdatavalid :  STD_LOGIC;
                signal ddr_sdram_s1_resetrequest_n :  STD_LOGIC;
                signal ddr_sdram_s1_resetrequest_n_from_sa :  STD_LOGIC;
                signal ddr_sdram_s1_waitrequest_n :  STD_LOGIC;
                signal ddr_sdram_s1_waitrequest_n_from_sa :  STD_LOGIC;
                signal ddr_sdram_s1_write :  STD_LOGIC;
                signal ddr_sdram_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_m1_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_m1_burstcount :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_m1_chipselect :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_debugaccess :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_endofpacket :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_latency_counter :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_read :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1_shift_register :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_m1_readdatavalid :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_waitrequest :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_write :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_m1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_arbiterlock :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_arbiterlock2 :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_burstcount :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_chipselect :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_debugaccess :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_endofpacket :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_read :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal flash_ssram_pipeline_bridge_s1_readdatavalid :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_reset_n :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_waitrequest :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_write :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal gpib_edm1_clock_0_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_0_in_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_edm1_clock_0_in_endofpacket :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal gpib_edm1_clock_0_in_read :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_0_in_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_0_in_reset_n :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_waitrequest :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_write :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_0_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_0_out_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_edm1_clock_0_out_endofpacket :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_granted_pll_s1 :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal gpib_edm1_clock_0_out_qualified_request_pll_s1 :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_read :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_read_data_valid_pll_s1 :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_0_out_requests_pll_s1 :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_reset_n :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_waitrequest :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_write :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_1_in_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpib_edm1_clock_1_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_1_in_endofpacket :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_endofpacket_from_sa :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_nativeaddress :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal gpib_edm1_clock_1_in_read :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal gpib_edm1_clock_1_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal gpib_edm1_clock_1_in_reset_n :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_waitrequest :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_waitrequest_from_sa :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_write :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal gpib_edm1_clock_1_out_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpib_edm1_clock_1_out_address_to_slave :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpib_edm1_clock_1_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_1_out_endofpacket :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_nativeaddress :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_read :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1 :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_reset_n :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_waitrequest :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_write :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal gpib_edm1_clock_2_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_2_in_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_edm1_clock_2_in_endofpacket :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_endofpacket_from_sa :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal gpib_edm1_clock_2_in_read :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_2_in_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_2_in_reset_n :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_waitrequest :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_waitrequest_from_sa :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_write :  STD_LOGIC;
                signal gpib_edm1_clock_2_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_2_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_2_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_2_out_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_edm1_clock_2_out_endofpacket :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_granted_ad7928_spi_control_port :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_read :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_read_data_valid_ad7928_spi_control_port :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_2_out_requests_ad7928_spi_control_port :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_reset_n :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_waitrequest :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_write :  STD_LOGIC;
                signal gpib_edm1_clock_2_out_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_3_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_3_in_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_edm1_clock_3_in_endofpacket :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_endofpacket_from_sa :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal gpib_edm1_clock_3_in_read :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_3_in_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_3_in_reset_n :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_waitrequest :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_waitrequest_from_sa :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_write :  STD_LOGIC;
                signal gpib_edm1_clock_3_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_3_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_3_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal gpib_edm1_clock_3_out_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_edm1_clock_3_out_endofpacket :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_read :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_read_data_valid_dac_ad5308_spi_control_port :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_reset_n :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_waitrequest :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_write :  STD_LOGIC;
                signal gpib_edm1_clock_3_out_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal gpib_leds_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpib_leds_s1_chipselect :  STD_LOGIC;
                signal gpib_leds_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpib_leds_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpib_leds_s1_reset_n :  STD_LOGIC;
                signal gpib_leds_s1_write_n :  STD_LOGIC;
                signal gpib_leds_s1_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpio1_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal gpio1_s1_chipselect :  STD_LOGIC;
                signal gpio1_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpio1_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpio1_s1_reset_n :  STD_LOGIC;
                signal gpio1_s1_write_n :  STD_LOGIC;
                signal gpio1_s1_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpio2_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal gpio2_s1_chipselect :  STD_LOGIC;
                signal gpio2_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpio2_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gpio2_s1_reset_n :  STD_LOGIC;
                signal gpio2_s1_write_n :  STD_LOGIC;
                signal gpio2_s1_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal high_res_timer_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal high_res_timer_s1_chipselect :  STD_LOGIC;
                signal high_res_timer_s1_irq :  STD_LOGIC;
                signal high_res_timer_s1_irq_from_sa :  STD_LOGIC;
                signal high_res_timer_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal high_res_timer_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal high_res_timer_s1_reset_n :  STD_LOGIC;
                signal high_res_timer_s1_write_n :  STD_LOGIC;
                signal high_res_timer_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal incoming_flash_ssram_tristate_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal incoming_flash_ssram_tristate_data_with_Xs_converted_to_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_MOSI_from_the_ad7928 :  STD_LOGIC;
                signal internal_MOSI_from_the_dac_ad5308 :  STD_LOGIC;
                signal internal_SCLK_from_the_ad7928 :  STD_LOGIC;
                signal internal_SCLK_from_the_dac_ad5308 :  STD_LOGIC;
                signal internal_SS_n_from_the_ad7928 :  STD_LOGIC;
                signal internal_SS_n_from_the_dac_ad5308 :  STD_LOGIC;
                signal internal_adsc_n_to_the_ssram :  STD_LOGIC;
                signal internal_bw_n_to_the_ssram :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_bwe_n_to_the_ssram :  STD_LOGIC;
                signal internal_chipenable1_n_to_the_ssram :  STD_LOGIC;
                signal internal_cpu_clk :  STD_LOGIC;
                signal internal_ddr_sdram_phy_clk_out :  STD_LOGIC;
                signal internal_flash_ssram_tristate_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal internal_local_init_done_from_the_ddr_sdram :  STD_LOGIC;
                signal internal_local_refresh_ack_from_the_ddr_sdram :  STD_LOGIC;
                signal internal_local_wdata_req_from_the_ddr_sdram :  STD_LOGIC;
                signal internal_mem_addr_from_the_ddr_sdram :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal internal_mem_ba_from_the_ddr_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_mem_cas_n_from_the_ddr_sdram :  STD_LOGIC;
                signal internal_mem_cke_from_the_ddr_sdram :  STD_LOGIC;
                signal internal_mem_cs_n_from_the_ddr_sdram :  STD_LOGIC;
                signal internal_mem_dm_from_the_ddr_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_mem_ras_n_from_the_ddr_sdram :  STD_LOGIC;
                signal internal_mem_we_n_from_the_ddr_sdram :  STD_LOGIC;
                signal internal_out_port_from_the_gpib_leds :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_out_port_from_the_gpio2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_out_port_from_the_led_pio :  STD_LOGIC;
                signal internal_outputenable_n_to_the_ssram :  STD_LOGIC;
                signal internal_pll_c2_out :  STD_LOGIC;
                signal internal_pll_c3_out :  STD_LOGIC;
                signal internal_read_n_to_the_cfi_flash :  STD_LOGIC;
                signal internal_reset_n_to_the_ssram :  STD_LOGIC;
                signal internal_reset_phy_clk_n_from_the_ddr_sdram :  STD_LOGIC;
                signal internal_select_n_to_the_cfi_flash :  STD_LOGIC;
                signal internal_write_n_to_the_cfi_flash :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_address :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_chipselect :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_read_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readyfordata :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reset_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_write_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal led_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal led_pio_s1_chipselect :  STD_LOGIC;
                signal led_pio_s1_readdata :  STD_LOGIC;
                signal led_pio_s1_readdata_from_sa :  STD_LOGIC;
                signal led_pio_s1_reset_n :  STD_LOGIC;
                signal led_pio_s1_write_n :  STD_LOGIC;
                signal led_pio_s1_writedata :  STD_LOGIC;
                signal module_input15 :  STD_LOGIC;
                signal module_input25 :  STD_LOGIC;
                signal module_input26 :  STD_LOGIC;
                signal module_input27 :  STD_LOGIC;
                signal module_input28 :  STD_LOGIC;
                signal onchip_memory_s1_address :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal onchip_memory_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal onchip_memory_s1_chipselect :  STD_LOGIC;
                signal onchip_memory_s1_clken :  STD_LOGIC;
                signal onchip_memory_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal onchip_memory_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal onchip_memory_s1_reset :  STD_LOGIC;
                signal onchip_memory_s1_write :  STD_LOGIC;
                signal onchip_memory_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal out_clk_ddr_sdram_aux_full_rate_clk :  STD_LOGIC;
                signal out_clk_ddr_sdram_aux_half_rate_clk :  STD_LOGIC;
                signal out_clk_ddr_sdram_phy_clk :  STD_LOGIC;
                signal out_clk_pll_c0 :  STD_LOGIC;
                signal out_clk_pll_c1 :  STD_LOGIC;
                signal out_clk_pll_c2 :  STD_LOGIC;
                signal out_clk_pll_c3 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_burstcount :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_chipselect :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_dbs_write_16 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_debugaccess :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_endofpacket :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_granted_ssram_s1 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_read :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pipeline_bridge_before_tristate_m1_readdatavalid :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_requests_ssram_s1 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_waitrequest :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_write :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pipeline_bridge_before_tristate_s1_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal pipeline_bridge_before_tristate_s1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_burstcount :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pipeline_bridge_before_tristate_s1_chipselect :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_debugaccess :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_endofpacket :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_endofpacket_from_sa :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal pipeline_bridge_before_tristate_s1_read :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pipeline_bridge_before_tristate_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pipeline_bridge_before_tristate_s1_readdatavalid :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_reset_n :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_waitrequest :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_waitrequest_from_sa :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_write :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pll_c2_out_reset_n :  STD_LOGIC;
                signal pll_c3_out_reset_n :  STD_LOGIC;
                signal pll_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pll_s1_chipselect :  STD_LOGIC;
                signal pll_s1_read :  STD_LOGIC;
                signal pll_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pll_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pll_s1_reset_n :  STD_LOGIC;
                signal pll_s1_resetrequest :  STD_LOGIC;
                signal pll_s1_resetrequest_from_sa :  STD_LOGIC;
                signal pll_s1_write :  STD_LOGIC;
                signal pll_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal registered_cpu_0_data_master_read_data_valid_onchip_memory_s1 :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_address :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal remote_update_cycloneiii_1_s1_chipselect :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_read :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal remote_update_cycloneiii_1_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal remote_update_cycloneiii_1_s1_reset :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_waitrequest :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_waitrequest_from_sa :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_write :  STD_LOGIC;
                signal remote_update_cycloneiii_1_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal reset_n_sources :  STD_LOGIC;
                signal sys_clk_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sys_clk_s1_chipselect :  STD_LOGIC;
                signal sys_clk_s1_irq :  STD_LOGIC;
                signal sys_clk_s1_irq_from_sa :  STD_LOGIC;
                signal sys_clk_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sys_clk_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sys_clk_s1_reset_n :  STD_LOGIC;
                signal sys_clk_s1_write_n :  STD_LOGIC;
                signal sys_clk_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);

begin

  --the_ad7928_spi_control_port, which is an e_instance
  the_ad7928_spi_control_port : ad7928_spi_control_port_arbitrator
    port map(
      ad7928_spi_control_port_address => ad7928_spi_control_port_address,
      ad7928_spi_control_port_chipselect => ad7928_spi_control_port_chipselect,
      ad7928_spi_control_port_dataavailable_from_sa => ad7928_spi_control_port_dataavailable_from_sa,
      ad7928_spi_control_port_endofpacket_from_sa => ad7928_spi_control_port_endofpacket_from_sa,
      ad7928_spi_control_port_irq_from_sa => ad7928_spi_control_port_irq_from_sa,
      ad7928_spi_control_port_read_n => ad7928_spi_control_port_read_n,
      ad7928_spi_control_port_readdata_from_sa => ad7928_spi_control_port_readdata_from_sa,
      ad7928_spi_control_port_readyfordata_from_sa => ad7928_spi_control_port_readyfordata_from_sa,
      ad7928_spi_control_port_reset_n => ad7928_spi_control_port_reset_n,
      ad7928_spi_control_port_write_n => ad7928_spi_control_port_write_n,
      ad7928_spi_control_port_writedata => ad7928_spi_control_port_writedata,
      d1_ad7928_spi_control_port_end_xfer => d1_ad7928_spi_control_port_end_xfer,
      gpib_edm1_clock_2_out_granted_ad7928_spi_control_port => gpib_edm1_clock_2_out_granted_ad7928_spi_control_port,
      gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port => gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port,
      gpib_edm1_clock_2_out_read_data_valid_ad7928_spi_control_port => gpib_edm1_clock_2_out_read_data_valid_ad7928_spi_control_port,
      gpib_edm1_clock_2_out_requests_ad7928_spi_control_port => gpib_edm1_clock_2_out_requests_ad7928_spi_control_port,
      ad7928_spi_control_port_dataavailable => ad7928_spi_control_port_dataavailable,
      ad7928_spi_control_port_endofpacket => ad7928_spi_control_port_endofpacket,
      ad7928_spi_control_port_irq => ad7928_spi_control_port_irq,
      ad7928_spi_control_port_readdata => ad7928_spi_control_port_readdata,
      ad7928_spi_control_port_readyfordata => ad7928_spi_control_port_readyfordata,
      clk => internal_cpu_clk,
      gpib_edm1_clock_2_out_address_to_slave => gpib_edm1_clock_2_out_address_to_slave,
      gpib_edm1_clock_2_out_nativeaddress => gpib_edm1_clock_2_out_nativeaddress,
      gpib_edm1_clock_2_out_read => gpib_edm1_clock_2_out_read,
      gpib_edm1_clock_2_out_write => gpib_edm1_clock_2_out_write,
      gpib_edm1_clock_2_out_writedata => gpib_edm1_clock_2_out_writedata,
      reset_n => cpu_clk_reset_n
    );


  --the_ad7928, which is an e_ptf_instance
  the_ad7928 : ad7928
    port map(
      MOSI => internal_MOSI_from_the_ad7928,
      SCLK => internal_SCLK_from_the_ad7928,
      SS_n => internal_SS_n_from_the_ad7928,
      data_to_cpu => ad7928_spi_control_port_readdata,
      dataavailable => ad7928_spi_control_port_dataavailable,
      endofpacket => ad7928_spi_control_port_endofpacket,
      irq => ad7928_spi_control_port_irq,
      readyfordata => ad7928_spi_control_port_readyfordata,
      MISO => MISO_to_the_ad7928,
      clk => internal_cpu_clk,
      data_from_cpu => ad7928_spi_control_port_writedata,
      mem_addr => ad7928_spi_control_port_address,
      read_n => ad7928_spi_control_port_read_n,
      reset_n => ad7928_spi_control_port_reset_n,
      spi_select => ad7928_spi_control_port_chipselect,
      write_n => ad7928_spi_control_port_write_n
    );


  --the_clock_crossing_0_s1, which is an e_instance
  the_clock_crossing_0_s1 : clock_crossing_0_s1_arbitrator
    port map(
      clock_crossing_0_s1_address => clock_crossing_0_s1_address,
      clock_crossing_0_s1_byteenable => clock_crossing_0_s1_byteenable,
      clock_crossing_0_s1_endofpacket_from_sa => clock_crossing_0_s1_endofpacket_from_sa,
      clock_crossing_0_s1_nativeaddress => clock_crossing_0_s1_nativeaddress,
      clock_crossing_0_s1_read => clock_crossing_0_s1_read,
      clock_crossing_0_s1_readdata_from_sa => clock_crossing_0_s1_readdata_from_sa,
      clock_crossing_0_s1_reset_n => clock_crossing_0_s1_reset_n,
      clock_crossing_0_s1_waitrequest_from_sa => clock_crossing_0_s1_waitrequest_from_sa,
      clock_crossing_0_s1_write => clock_crossing_0_s1_write,
      clock_crossing_0_s1_writedata => clock_crossing_0_s1_writedata,
      cpu_0_data_master_granted_clock_crossing_0_s1 => cpu_0_data_master_granted_clock_crossing_0_s1,
      cpu_0_data_master_qualified_request_clock_crossing_0_s1 => cpu_0_data_master_qualified_request_clock_crossing_0_s1,
      cpu_0_data_master_read_data_valid_clock_crossing_0_s1 => cpu_0_data_master_read_data_valid_clock_crossing_0_s1,
      cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register => cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register,
      cpu_0_data_master_requests_clock_crossing_0_s1 => cpu_0_data_master_requests_clock_crossing_0_s1,
      cpu_0_instruction_master_granted_clock_crossing_0_s1 => cpu_0_instruction_master_granted_clock_crossing_0_s1,
      cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 => cpu_0_instruction_master_qualified_request_clock_crossing_0_s1,
      cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1 => cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1,
      cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register => cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register,
      cpu_0_instruction_master_requests_clock_crossing_0_s1 => cpu_0_instruction_master_requests_clock_crossing_0_s1,
      d1_clock_crossing_0_s1_end_xfer => d1_clock_crossing_0_s1_end_xfer,
      clk => internal_cpu_clk,
      clock_crossing_0_s1_endofpacket => clock_crossing_0_s1_endofpacket,
      clock_crossing_0_s1_readdata => clock_crossing_0_s1_readdata,
      clock_crossing_0_s1_readdatavalid => clock_crossing_0_s1_readdatavalid,
      clock_crossing_0_s1_waitrequest => clock_crossing_0_s1_waitrequest,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_waitrequest => cpu_0_data_master_waitrequest,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      cpu_0_instruction_master_address_to_slave => cpu_0_instruction_master_address_to_slave,
      cpu_0_instruction_master_read => cpu_0_instruction_master_read,
      reset_n => cpu_clk_reset_n
    );


  --the_clock_crossing_0_m1, which is an e_instance
  the_clock_crossing_0_m1 : clock_crossing_0_m1_arbitrator
    port map(
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_endofpacket => clock_crossing_0_m1_endofpacket,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_readdata => clock_crossing_0_m1_readdata,
      clock_crossing_0_m1_readdatavalid => clock_crossing_0_m1_readdatavalid,
      clock_crossing_0_m1_reset_n => clock_crossing_0_m1_reset_n,
      clock_crossing_0_m1_waitrequest => clock_crossing_0_m1_waitrequest,
      clk => internal_pll_c2_out,
      clock_crossing_0_m1_address => clock_crossing_0_m1_address,
      clock_crossing_0_m1_byteenable => clock_crossing_0_m1_byteenable,
      clock_crossing_0_m1_granted_gpib_edm1_clock_2_in => clock_crossing_0_m1_granted_gpib_edm1_clock_2_in,
      clock_crossing_0_m1_granted_gpib_edm1_clock_3_in => clock_crossing_0_m1_granted_gpib_edm1_clock_3_in,
      clock_crossing_0_m1_granted_gpib_leds_s1 => clock_crossing_0_m1_granted_gpib_leds_s1,
      clock_crossing_0_m1_granted_gpio1_s1 => clock_crossing_0_m1_granted_gpio1_s1,
      clock_crossing_0_m1_granted_gpio2_s1 => clock_crossing_0_m1_granted_gpio2_s1,
      clock_crossing_0_m1_granted_high_res_timer_s1 => clock_crossing_0_m1_granted_high_res_timer_s1,
      clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave => clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave,
      clock_crossing_0_m1_granted_led_pio_s1 => clock_crossing_0_m1_granted_led_pio_s1,
      clock_crossing_0_m1_granted_sys_clk_s1 => clock_crossing_0_m1_granted_sys_clk_s1,
      clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in => clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in,
      clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in => clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in,
      clock_crossing_0_m1_qualified_request_gpib_leds_s1 => clock_crossing_0_m1_qualified_request_gpib_leds_s1,
      clock_crossing_0_m1_qualified_request_gpio1_s1 => clock_crossing_0_m1_qualified_request_gpio1_s1,
      clock_crossing_0_m1_qualified_request_gpio2_s1 => clock_crossing_0_m1_qualified_request_gpio2_s1,
      clock_crossing_0_m1_qualified_request_high_res_timer_s1 => clock_crossing_0_m1_qualified_request_high_res_timer_s1,
      clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave => clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave,
      clock_crossing_0_m1_qualified_request_led_pio_s1 => clock_crossing_0_m1_qualified_request_led_pio_s1,
      clock_crossing_0_m1_qualified_request_sys_clk_s1 => clock_crossing_0_m1_qualified_request_sys_clk_s1,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in => clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in,
      clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in => clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in,
      clock_crossing_0_m1_read_data_valid_gpib_leds_s1 => clock_crossing_0_m1_read_data_valid_gpib_leds_s1,
      clock_crossing_0_m1_read_data_valid_gpio1_s1 => clock_crossing_0_m1_read_data_valid_gpio1_s1,
      clock_crossing_0_m1_read_data_valid_gpio2_s1 => clock_crossing_0_m1_read_data_valid_gpio2_s1,
      clock_crossing_0_m1_read_data_valid_high_res_timer_s1 => clock_crossing_0_m1_read_data_valid_high_res_timer_s1,
      clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave => clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
      clock_crossing_0_m1_read_data_valid_led_pio_s1 => clock_crossing_0_m1_read_data_valid_led_pio_s1,
      clock_crossing_0_m1_read_data_valid_sys_clk_s1 => clock_crossing_0_m1_read_data_valid_sys_clk_s1,
      clock_crossing_0_m1_requests_gpib_edm1_clock_2_in => clock_crossing_0_m1_requests_gpib_edm1_clock_2_in,
      clock_crossing_0_m1_requests_gpib_edm1_clock_3_in => clock_crossing_0_m1_requests_gpib_edm1_clock_3_in,
      clock_crossing_0_m1_requests_gpib_leds_s1 => clock_crossing_0_m1_requests_gpib_leds_s1,
      clock_crossing_0_m1_requests_gpio1_s1 => clock_crossing_0_m1_requests_gpio1_s1,
      clock_crossing_0_m1_requests_gpio2_s1 => clock_crossing_0_m1_requests_gpio2_s1,
      clock_crossing_0_m1_requests_high_res_timer_s1 => clock_crossing_0_m1_requests_high_res_timer_s1,
      clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave => clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave,
      clock_crossing_0_m1_requests_led_pio_s1 => clock_crossing_0_m1_requests_led_pio_s1,
      clock_crossing_0_m1_requests_sys_clk_s1 => clock_crossing_0_m1_requests_sys_clk_s1,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      d1_gpib_edm1_clock_2_in_end_xfer => d1_gpib_edm1_clock_2_in_end_xfer,
      d1_gpib_edm1_clock_3_in_end_xfer => d1_gpib_edm1_clock_3_in_end_xfer,
      d1_gpib_leds_s1_end_xfer => d1_gpib_leds_s1_end_xfer,
      d1_gpio1_s1_end_xfer => d1_gpio1_s1_end_xfer,
      d1_gpio2_s1_end_xfer => d1_gpio2_s1_end_xfer,
      d1_high_res_timer_s1_end_xfer => d1_high_res_timer_s1_end_xfer,
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      d1_led_pio_s1_end_xfer => d1_led_pio_s1_end_xfer,
      d1_sys_clk_s1_end_xfer => d1_sys_clk_s1_end_xfer,
      gpib_edm1_clock_2_in_endofpacket_from_sa => gpib_edm1_clock_2_in_endofpacket_from_sa,
      gpib_edm1_clock_2_in_readdata_from_sa => gpib_edm1_clock_2_in_readdata_from_sa,
      gpib_edm1_clock_2_in_waitrequest_from_sa => gpib_edm1_clock_2_in_waitrequest_from_sa,
      gpib_edm1_clock_3_in_endofpacket_from_sa => gpib_edm1_clock_3_in_endofpacket_from_sa,
      gpib_edm1_clock_3_in_readdata_from_sa => gpib_edm1_clock_3_in_readdata_from_sa,
      gpib_edm1_clock_3_in_waitrequest_from_sa => gpib_edm1_clock_3_in_waitrequest_from_sa,
      gpib_leds_s1_readdata_from_sa => gpib_leds_s1_readdata_from_sa,
      gpio1_s1_readdata_from_sa => gpio1_s1_readdata_from_sa,
      gpio2_s1_readdata_from_sa => gpio2_s1_readdata_from_sa,
      high_res_timer_s1_readdata_from_sa => high_res_timer_s1_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      led_pio_s1_readdata_from_sa => led_pio_s1_readdata_from_sa,
      reset_n => pll_c2_out_reset_n,
      sys_clk_s1_readdata_from_sa => sys_clk_s1_readdata_from_sa
    );


  --the_clock_crossing_0, which is an e_ptf_instance
  the_clock_crossing_0 : clock_crossing_0
    port map(
      master_address => clock_crossing_0_m1_address,
      master_byteenable => clock_crossing_0_m1_byteenable,
      master_nativeaddress => clock_crossing_0_m1_nativeaddress,
      master_read => clock_crossing_0_m1_read,
      master_write => clock_crossing_0_m1_write,
      master_writedata => clock_crossing_0_m1_writedata,
      slave_endofpacket => clock_crossing_0_s1_endofpacket,
      slave_readdata => clock_crossing_0_s1_readdata,
      slave_readdatavalid => clock_crossing_0_s1_readdatavalid,
      slave_waitrequest => clock_crossing_0_s1_waitrequest,
      master_clk => internal_pll_c2_out,
      master_endofpacket => clock_crossing_0_m1_endofpacket,
      master_readdata => clock_crossing_0_m1_readdata,
      master_readdatavalid => clock_crossing_0_m1_readdatavalid,
      master_reset_n => clock_crossing_0_m1_reset_n,
      master_waitrequest => clock_crossing_0_m1_waitrequest,
      slave_address => clock_crossing_0_s1_address,
      slave_byteenable => clock_crossing_0_s1_byteenable,
      slave_clk => internal_cpu_clk,
      slave_nativeaddress => clock_crossing_0_s1_nativeaddress,
      slave_read => clock_crossing_0_s1_read,
      slave_reset_n => clock_crossing_0_s1_reset_n,
      slave_write => clock_crossing_0_s1_write,
      slave_writedata => clock_crossing_0_s1_writedata
    );


  --the_cpu_0_jtag_debug_module, which is an e_instance
  the_cpu_0_jtag_debug_module : cpu_0_jtag_debug_module_arbitrator
    port map(
      cpu_0_data_master_granted_cpu_0_jtag_debug_module => cpu_0_data_master_granted_cpu_0_jtag_debug_module,
      cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module => cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module,
      cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module => cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module,
      cpu_0_data_master_requests_cpu_0_jtag_debug_module => cpu_0_data_master_requests_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_granted_cpu_0_jtag_debug_module => cpu_0_instruction_master_granted_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module => cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module => cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_requests_cpu_0_jtag_debug_module => cpu_0_instruction_master_requests_cpu_0_jtag_debug_module,
      cpu_0_jtag_debug_module_address => cpu_0_jtag_debug_module_address,
      cpu_0_jtag_debug_module_begintransfer => cpu_0_jtag_debug_module_begintransfer,
      cpu_0_jtag_debug_module_byteenable => cpu_0_jtag_debug_module_byteenable,
      cpu_0_jtag_debug_module_chipselect => cpu_0_jtag_debug_module_chipselect,
      cpu_0_jtag_debug_module_debugaccess => cpu_0_jtag_debug_module_debugaccess,
      cpu_0_jtag_debug_module_readdata_from_sa => cpu_0_jtag_debug_module_readdata_from_sa,
      cpu_0_jtag_debug_module_reset_n => cpu_0_jtag_debug_module_reset_n,
      cpu_0_jtag_debug_module_resetrequest_from_sa => cpu_0_jtag_debug_module_resetrequest_from_sa,
      cpu_0_jtag_debug_module_write => cpu_0_jtag_debug_module_write,
      cpu_0_jtag_debug_module_writedata => cpu_0_jtag_debug_module_writedata,
      d1_cpu_0_jtag_debug_module_end_xfer => d1_cpu_0_jtag_debug_module_end_xfer,
      clk => internal_cpu_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_debugaccess => cpu_0_data_master_debugaccess,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_waitrequest => cpu_0_data_master_waitrequest,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      cpu_0_instruction_master_address_to_slave => cpu_0_instruction_master_address_to_slave,
      cpu_0_instruction_master_read => cpu_0_instruction_master_read,
      cpu_0_jtag_debug_module_readdata => cpu_0_jtag_debug_module_readdata,
      cpu_0_jtag_debug_module_resetrequest => cpu_0_jtag_debug_module_resetrequest,
      reset_n => cpu_clk_reset_n
    );


  --the_cpu_0_data_master, which is an e_instance
  the_cpu_0_data_master : cpu_0_data_master_arbitrator
    port map(
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_irq => cpu_0_data_master_irq,
      cpu_0_data_master_readdata => cpu_0_data_master_readdata,
      cpu_0_data_master_waitrequest => cpu_0_data_master_waitrequest,
      ad7928_spi_control_port_irq_from_sa => ad7928_spi_control_port_irq_from_sa,
      clk => internal_cpu_clk,
      clock_crossing_0_s1_readdata_from_sa => clock_crossing_0_s1_readdata_from_sa,
      clock_crossing_0_s1_waitrequest_from_sa => clock_crossing_0_s1_waitrequest_from_sa,
      cpu_0_data_master_address => cpu_0_data_master_address,
      cpu_0_data_master_granted_clock_crossing_0_s1 => cpu_0_data_master_granted_clock_crossing_0_s1,
      cpu_0_data_master_granted_cpu_0_jtag_debug_module => cpu_0_data_master_granted_cpu_0_jtag_debug_module,
      cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 => cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1,
      cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 => cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1,
      cpu_0_data_master_granted_gpib_edm1_clock_0_in => cpu_0_data_master_granted_gpib_edm1_clock_0_in,
      cpu_0_data_master_granted_gpib_edm1_clock_1_in => cpu_0_data_master_granted_gpib_edm1_clock_1_in,
      cpu_0_data_master_granted_onchip_memory_s1 => cpu_0_data_master_granted_onchip_memory_s1,
      cpu_0_data_master_qualified_request_clock_crossing_0_s1 => cpu_0_data_master_qualified_request_clock_crossing_0_s1,
      cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module => cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module,
      cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 => cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1,
      cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 => cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1,
      cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in => cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in,
      cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in => cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in,
      cpu_0_data_master_qualified_request_onchip_memory_s1 => cpu_0_data_master_qualified_request_onchip_memory_s1,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_read_data_valid_clock_crossing_0_s1 => cpu_0_data_master_read_data_valid_clock_crossing_0_s1,
      cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register => cpu_0_data_master_read_data_valid_clock_crossing_0_s1_shift_register,
      cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module => cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module,
      cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 => cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1,
      cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register => cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
      cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1 => cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1,
      cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register => cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
      cpu_0_data_master_read_data_valid_gpib_edm1_clock_0_in => cpu_0_data_master_read_data_valid_gpib_edm1_clock_0_in,
      cpu_0_data_master_read_data_valid_gpib_edm1_clock_1_in => cpu_0_data_master_read_data_valid_gpib_edm1_clock_1_in,
      cpu_0_data_master_read_data_valid_onchip_memory_s1 => cpu_0_data_master_read_data_valid_onchip_memory_s1,
      cpu_0_data_master_requests_clock_crossing_0_s1 => cpu_0_data_master_requests_clock_crossing_0_s1,
      cpu_0_data_master_requests_cpu_0_jtag_debug_module => cpu_0_data_master_requests_cpu_0_jtag_debug_module,
      cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 => cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1,
      cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 => cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1,
      cpu_0_data_master_requests_gpib_edm1_clock_0_in => cpu_0_data_master_requests_gpib_edm1_clock_0_in,
      cpu_0_data_master_requests_gpib_edm1_clock_1_in => cpu_0_data_master_requests_gpib_edm1_clock_1_in,
      cpu_0_data_master_requests_onchip_memory_s1 => cpu_0_data_master_requests_onchip_memory_s1,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_jtag_debug_module_readdata_from_sa => cpu_0_jtag_debug_module_readdata_from_sa,
      cpu_clk => internal_cpu_clk,
      cpu_clk_reset_n => cpu_clk_reset_n,
      cpu_ddr_clock_bridge_s1_readdata_from_sa => cpu_ddr_clock_bridge_s1_readdata_from_sa,
      cpu_ddr_clock_bridge_s1_waitrequest_from_sa => cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
      d1_clock_crossing_0_s1_end_xfer => d1_clock_crossing_0_s1_end_xfer,
      d1_cpu_0_jtag_debug_module_end_xfer => d1_cpu_0_jtag_debug_module_end_xfer,
      d1_cpu_ddr_clock_bridge_s1_end_xfer => d1_cpu_ddr_clock_bridge_s1_end_xfer,
      d1_flash_ssram_pipeline_bridge_s1_end_xfer => d1_flash_ssram_pipeline_bridge_s1_end_xfer,
      d1_gpib_edm1_clock_0_in_end_xfer => d1_gpib_edm1_clock_0_in_end_xfer,
      d1_gpib_edm1_clock_1_in_end_xfer => d1_gpib_edm1_clock_1_in_end_xfer,
      d1_onchip_memory_s1_end_xfer => d1_onchip_memory_s1_end_xfer,
      dac_ad5308_spi_control_port_irq_from_sa => dac_ad5308_spi_control_port_irq_from_sa,
      flash_ssram_pipeline_bridge_s1_readdata_from_sa => flash_ssram_pipeline_bridge_s1_readdata_from_sa,
      flash_ssram_pipeline_bridge_s1_waitrequest_from_sa => flash_ssram_pipeline_bridge_s1_waitrequest_from_sa,
      gpib_edm1_clock_0_in_readdata_from_sa => gpib_edm1_clock_0_in_readdata_from_sa,
      gpib_edm1_clock_0_in_waitrequest_from_sa => gpib_edm1_clock_0_in_waitrequest_from_sa,
      gpib_edm1_clock_1_in_readdata_from_sa => gpib_edm1_clock_1_in_readdata_from_sa,
      gpib_edm1_clock_1_in_waitrequest_from_sa => gpib_edm1_clock_1_in_waitrequest_from_sa,
      high_res_timer_s1_irq_from_sa => high_res_timer_s1_irq_from_sa,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      onchip_memory_s1_readdata_from_sa => onchip_memory_s1_readdata_from_sa,
      registered_cpu_0_data_master_read_data_valid_onchip_memory_s1 => registered_cpu_0_data_master_read_data_valid_onchip_memory_s1,
      reset_n => cpu_clk_reset_n,
      sys_clk_s1_irq_from_sa => sys_clk_s1_irq_from_sa
    );


  --the_cpu_0_instruction_master, which is an e_instance
  the_cpu_0_instruction_master : cpu_0_instruction_master_arbitrator
    port map(
      cpu_0_instruction_master_address_to_slave => cpu_0_instruction_master_address_to_slave,
      cpu_0_instruction_master_readdata => cpu_0_instruction_master_readdata,
      cpu_0_instruction_master_waitrequest => cpu_0_instruction_master_waitrequest,
      clk => internal_cpu_clk,
      clock_crossing_0_s1_readdata_from_sa => clock_crossing_0_s1_readdata_from_sa,
      clock_crossing_0_s1_waitrequest_from_sa => clock_crossing_0_s1_waitrequest_from_sa,
      cpu_0_instruction_master_address => cpu_0_instruction_master_address,
      cpu_0_instruction_master_granted_clock_crossing_0_s1 => cpu_0_instruction_master_granted_clock_crossing_0_s1,
      cpu_0_instruction_master_granted_cpu_0_jtag_debug_module => cpu_0_instruction_master_granted_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 => cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1,
      cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 => cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1,
      cpu_0_instruction_master_granted_onchip_memory_s1 => cpu_0_instruction_master_granted_onchip_memory_s1,
      cpu_0_instruction_master_qualified_request_clock_crossing_0_s1 => cpu_0_instruction_master_qualified_request_clock_crossing_0_s1,
      cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module => cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 => cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1,
      cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 => cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1,
      cpu_0_instruction_master_qualified_request_onchip_memory_s1 => cpu_0_instruction_master_qualified_request_onchip_memory_s1,
      cpu_0_instruction_master_read => cpu_0_instruction_master_read,
      cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1 => cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1,
      cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register => cpu_0_instruction_master_read_data_valid_clock_crossing_0_s1_shift_register,
      cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module => cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 => cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1,
      cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register => cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
      cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1 => cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1,
      cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register => cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
      cpu_0_instruction_master_read_data_valid_onchip_memory_s1 => cpu_0_instruction_master_read_data_valid_onchip_memory_s1,
      cpu_0_instruction_master_requests_clock_crossing_0_s1 => cpu_0_instruction_master_requests_clock_crossing_0_s1,
      cpu_0_instruction_master_requests_cpu_0_jtag_debug_module => cpu_0_instruction_master_requests_cpu_0_jtag_debug_module,
      cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 => cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1,
      cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 => cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1,
      cpu_0_instruction_master_requests_onchip_memory_s1 => cpu_0_instruction_master_requests_onchip_memory_s1,
      cpu_0_jtag_debug_module_readdata_from_sa => cpu_0_jtag_debug_module_readdata_from_sa,
      cpu_ddr_clock_bridge_s1_readdata_from_sa => cpu_ddr_clock_bridge_s1_readdata_from_sa,
      cpu_ddr_clock_bridge_s1_waitrequest_from_sa => cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
      d1_clock_crossing_0_s1_end_xfer => d1_clock_crossing_0_s1_end_xfer,
      d1_cpu_0_jtag_debug_module_end_xfer => d1_cpu_0_jtag_debug_module_end_xfer,
      d1_cpu_ddr_clock_bridge_s1_end_xfer => d1_cpu_ddr_clock_bridge_s1_end_xfer,
      d1_flash_ssram_pipeline_bridge_s1_end_xfer => d1_flash_ssram_pipeline_bridge_s1_end_xfer,
      d1_onchip_memory_s1_end_xfer => d1_onchip_memory_s1_end_xfer,
      flash_ssram_pipeline_bridge_s1_readdata_from_sa => flash_ssram_pipeline_bridge_s1_readdata_from_sa,
      flash_ssram_pipeline_bridge_s1_waitrequest_from_sa => flash_ssram_pipeline_bridge_s1_waitrequest_from_sa,
      onchip_memory_s1_readdata_from_sa => onchip_memory_s1_readdata_from_sa,
      reset_n => cpu_clk_reset_n
    );


  --the_cpu_0, which is an e_ptf_instance
  the_cpu_0 : cpu_0
    port map(
      d_address => cpu_0_data_master_address,
      d_byteenable => cpu_0_data_master_byteenable,
      d_read => cpu_0_data_master_read,
      d_write => cpu_0_data_master_write,
      d_writedata => cpu_0_data_master_writedata,
      i_address => cpu_0_instruction_master_address,
      i_read => cpu_0_instruction_master_read,
      jtag_debug_module_debugaccess_to_roms => cpu_0_data_master_debugaccess,
      jtag_debug_module_readdata => cpu_0_jtag_debug_module_readdata,
      jtag_debug_module_resetrequest => cpu_0_jtag_debug_module_resetrequest,
      clk => internal_cpu_clk,
      d_irq => cpu_0_data_master_irq,
      d_readdata => cpu_0_data_master_readdata,
      d_waitrequest => cpu_0_data_master_waitrequest,
      i_readdata => cpu_0_instruction_master_readdata,
      i_waitrequest => cpu_0_instruction_master_waitrequest,
      jtag_debug_module_address => cpu_0_jtag_debug_module_address,
      jtag_debug_module_begintransfer => cpu_0_jtag_debug_module_begintransfer,
      jtag_debug_module_byteenable => cpu_0_jtag_debug_module_byteenable,
      jtag_debug_module_debugaccess => cpu_0_jtag_debug_module_debugaccess,
      jtag_debug_module_select => cpu_0_jtag_debug_module_chipselect,
      jtag_debug_module_write => cpu_0_jtag_debug_module_write,
      jtag_debug_module_writedata => cpu_0_jtag_debug_module_writedata,
      reset_n => cpu_0_jtag_debug_module_reset_n
    );


  --the_cpu_ddr_clock_bridge_s1, which is an e_instance
  the_cpu_ddr_clock_bridge_s1 : cpu_ddr_clock_bridge_s1_arbitrator
    port map(
      cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1 => cpu_0_data_master_granted_cpu_ddr_clock_bridge_s1,
      cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1 => cpu_0_data_master_qualified_request_cpu_ddr_clock_bridge_s1,
      cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 => cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1,
      cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register => cpu_0_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
      cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1 => cpu_0_data_master_requests_cpu_ddr_clock_bridge_s1,
      cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1 => cpu_0_instruction_master_granted_cpu_ddr_clock_bridge_s1,
      cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 => cpu_0_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1,
      cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 => cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1,
      cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register => cpu_0_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
      cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1 => cpu_0_instruction_master_requests_cpu_ddr_clock_bridge_s1,
      cpu_ddr_clock_bridge_s1_address => cpu_ddr_clock_bridge_s1_address,
      cpu_ddr_clock_bridge_s1_byteenable => cpu_ddr_clock_bridge_s1_byteenable,
      cpu_ddr_clock_bridge_s1_endofpacket_from_sa => cpu_ddr_clock_bridge_s1_endofpacket_from_sa,
      cpu_ddr_clock_bridge_s1_nativeaddress => cpu_ddr_clock_bridge_s1_nativeaddress,
      cpu_ddr_clock_bridge_s1_read => cpu_ddr_clock_bridge_s1_read,
      cpu_ddr_clock_bridge_s1_readdata_from_sa => cpu_ddr_clock_bridge_s1_readdata_from_sa,
      cpu_ddr_clock_bridge_s1_reset_n => cpu_ddr_clock_bridge_s1_reset_n,
      cpu_ddr_clock_bridge_s1_waitrequest_from_sa => cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
      cpu_ddr_clock_bridge_s1_write => cpu_ddr_clock_bridge_s1_write,
      cpu_ddr_clock_bridge_s1_writedata => cpu_ddr_clock_bridge_s1_writedata,
      d1_cpu_ddr_clock_bridge_s1_end_xfer => d1_cpu_ddr_clock_bridge_s1_end_xfer,
      clk => internal_cpu_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_waitrequest => cpu_0_data_master_waitrequest,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      cpu_0_instruction_master_address_to_slave => cpu_0_instruction_master_address_to_slave,
      cpu_0_instruction_master_read => cpu_0_instruction_master_read,
      cpu_ddr_clock_bridge_s1_endofpacket => cpu_ddr_clock_bridge_s1_endofpacket,
      cpu_ddr_clock_bridge_s1_readdata => cpu_ddr_clock_bridge_s1_readdata,
      cpu_ddr_clock_bridge_s1_readdatavalid => cpu_ddr_clock_bridge_s1_readdatavalid,
      cpu_ddr_clock_bridge_s1_waitrequest => cpu_ddr_clock_bridge_s1_waitrequest,
      reset_n => cpu_clk_reset_n
    );


  --the_cpu_ddr_clock_bridge_m1, which is an e_instance
  the_cpu_ddr_clock_bridge_m1 : cpu_ddr_clock_bridge_m1_arbitrator
    port map(
      cpu_ddr_clock_bridge_m1_address_to_slave => cpu_ddr_clock_bridge_m1_address_to_slave,
      cpu_ddr_clock_bridge_m1_latency_counter => cpu_ddr_clock_bridge_m1_latency_counter,
      cpu_ddr_clock_bridge_m1_readdata => cpu_ddr_clock_bridge_m1_readdata,
      cpu_ddr_clock_bridge_m1_readdatavalid => cpu_ddr_clock_bridge_m1_readdatavalid,
      cpu_ddr_clock_bridge_m1_reset_n => cpu_ddr_clock_bridge_m1_reset_n,
      cpu_ddr_clock_bridge_m1_waitrequest => cpu_ddr_clock_bridge_m1_waitrequest,
      clk => internal_ddr_sdram_phy_clk_out,
      cpu_ddr_clock_bridge_m1_address => cpu_ddr_clock_bridge_m1_address,
      cpu_ddr_clock_bridge_m1_byteenable => cpu_ddr_clock_bridge_m1_byteenable,
      cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 => cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1,
      cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 => cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1,
      cpu_ddr_clock_bridge_m1_read => cpu_ddr_clock_bridge_m1_read,
      cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1 => cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1,
      cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1_shift_register => cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1_shift_register,
      cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 => cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1,
      cpu_ddr_clock_bridge_m1_write => cpu_ddr_clock_bridge_m1_write,
      cpu_ddr_clock_bridge_m1_writedata => cpu_ddr_clock_bridge_m1_writedata,
      d1_ddr_sdram_s1_end_xfer => d1_ddr_sdram_s1_end_xfer,
      ddr_sdram_s1_readdata_from_sa => ddr_sdram_s1_readdata_from_sa,
      ddr_sdram_s1_waitrequest_n_from_sa => ddr_sdram_s1_waitrequest_n_from_sa,
      reset_n => ddr_sdram_phy_clk_out_reset_n
    );


  --the_cpu_ddr_clock_bridge, which is an e_ptf_instance
  the_cpu_ddr_clock_bridge : cpu_ddr_clock_bridge
    port map(
      master_address => cpu_ddr_clock_bridge_m1_address,
      master_byteenable => cpu_ddr_clock_bridge_m1_byteenable,
      master_nativeaddress => cpu_ddr_clock_bridge_m1_nativeaddress,
      master_read => cpu_ddr_clock_bridge_m1_read,
      master_write => cpu_ddr_clock_bridge_m1_write,
      master_writedata => cpu_ddr_clock_bridge_m1_writedata,
      slave_endofpacket => cpu_ddr_clock_bridge_s1_endofpacket,
      slave_readdata => cpu_ddr_clock_bridge_s1_readdata,
      slave_readdatavalid => cpu_ddr_clock_bridge_s1_readdatavalid,
      slave_waitrequest => cpu_ddr_clock_bridge_s1_waitrequest,
      master_clk => internal_ddr_sdram_phy_clk_out,
      master_endofpacket => cpu_ddr_clock_bridge_m1_endofpacket,
      master_readdata => cpu_ddr_clock_bridge_m1_readdata,
      master_readdatavalid => cpu_ddr_clock_bridge_m1_readdatavalid,
      master_reset_n => cpu_ddr_clock_bridge_m1_reset_n,
      master_waitrequest => cpu_ddr_clock_bridge_m1_waitrequest,
      slave_address => cpu_ddr_clock_bridge_s1_address,
      slave_byteenable => cpu_ddr_clock_bridge_s1_byteenable,
      slave_clk => internal_cpu_clk,
      slave_nativeaddress => cpu_ddr_clock_bridge_s1_nativeaddress,
      slave_read => cpu_ddr_clock_bridge_s1_read,
      slave_reset_n => cpu_ddr_clock_bridge_s1_reset_n,
      slave_write => cpu_ddr_clock_bridge_s1_write,
      slave_writedata => cpu_ddr_clock_bridge_s1_writedata
    );


  --the_dac_ad5308_spi_control_port, which is an e_instance
  the_dac_ad5308_spi_control_port : dac_ad5308_spi_control_port_arbitrator
    port map(
      d1_dac_ad5308_spi_control_port_end_xfer => d1_dac_ad5308_spi_control_port_end_xfer,
      dac_ad5308_spi_control_port_address => dac_ad5308_spi_control_port_address,
      dac_ad5308_spi_control_port_chipselect => dac_ad5308_spi_control_port_chipselect,
      dac_ad5308_spi_control_port_dataavailable_from_sa => dac_ad5308_spi_control_port_dataavailable_from_sa,
      dac_ad5308_spi_control_port_endofpacket_from_sa => dac_ad5308_spi_control_port_endofpacket_from_sa,
      dac_ad5308_spi_control_port_irq_from_sa => dac_ad5308_spi_control_port_irq_from_sa,
      dac_ad5308_spi_control_port_read_n => dac_ad5308_spi_control_port_read_n,
      dac_ad5308_spi_control_port_readdata_from_sa => dac_ad5308_spi_control_port_readdata_from_sa,
      dac_ad5308_spi_control_port_readyfordata_from_sa => dac_ad5308_spi_control_port_readyfordata_from_sa,
      dac_ad5308_spi_control_port_reset_n => dac_ad5308_spi_control_port_reset_n,
      dac_ad5308_spi_control_port_write_n => dac_ad5308_spi_control_port_write_n,
      dac_ad5308_spi_control_port_writedata => dac_ad5308_spi_control_port_writedata,
      gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port => gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port,
      gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port => gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port,
      gpib_edm1_clock_3_out_read_data_valid_dac_ad5308_spi_control_port => gpib_edm1_clock_3_out_read_data_valid_dac_ad5308_spi_control_port,
      gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port => gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port,
      clk => internal_cpu_clk,
      dac_ad5308_spi_control_port_dataavailable => dac_ad5308_spi_control_port_dataavailable,
      dac_ad5308_spi_control_port_endofpacket => dac_ad5308_spi_control_port_endofpacket,
      dac_ad5308_spi_control_port_irq => dac_ad5308_spi_control_port_irq,
      dac_ad5308_spi_control_port_readdata => dac_ad5308_spi_control_port_readdata,
      dac_ad5308_spi_control_port_readyfordata => dac_ad5308_spi_control_port_readyfordata,
      gpib_edm1_clock_3_out_address_to_slave => gpib_edm1_clock_3_out_address_to_slave,
      gpib_edm1_clock_3_out_nativeaddress => gpib_edm1_clock_3_out_nativeaddress,
      gpib_edm1_clock_3_out_read => gpib_edm1_clock_3_out_read,
      gpib_edm1_clock_3_out_write => gpib_edm1_clock_3_out_write,
      gpib_edm1_clock_3_out_writedata => gpib_edm1_clock_3_out_writedata,
      reset_n => cpu_clk_reset_n
    );


  --the_dac_ad5308, which is an e_ptf_instance
  the_dac_ad5308 : dac_ad5308
    port map(
      MOSI => internal_MOSI_from_the_dac_ad5308,
      SCLK => internal_SCLK_from_the_dac_ad5308,
      SS_n => internal_SS_n_from_the_dac_ad5308,
      data_to_cpu => dac_ad5308_spi_control_port_readdata,
      dataavailable => dac_ad5308_spi_control_port_dataavailable,
      endofpacket => dac_ad5308_spi_control_port_endofpacket,
      irq => dac_ad5308_spi_control_port_irq,
      readyfordata => dac_ad5308_spi_control_port_readyfordata,
      MISO => MISO_to_the_dac_ad5308,
      clk => internal_cpu_clk,
      data_from_cpu => dac_ad5308_spi_control_port_writedata,
      mem_addr => dac_ad5308_spi_control_port_address,
      read_n => dac_ad5308_spi_control_port_read_n,
      reset_n => dac_ad5308_spi_control_port_reset_n,
      spi_select => dac_ad5308_spi_control_port_chipselect,
      write_n => dac_ad5308_spi_control_port_write_n
    );


  --the_ddr_sdram_s1, which is an e_instance
  the_ddr_sdram_s1 : ddr_sdram_s1_arbitrator
    port map(
      cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1 => cpu_ddr_clock_bridge_m1_granted_ddr_sdram_s1,
      cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1 => cpu_ddr_clock_bridge_m1_qualified_request_ddr_sdram_s1,
      cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1 => cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1,
      cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1_shift_register => cpu_ddr_clock_bridge_m1_read_data_valid_ddr_sdram_s1_shift_register,
      cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1 => cpu_ddr_clock_bridge_m1_requests_ddr_sdram_s1,
      d1_ddr_sdram_s1_end_xfer => d1_ddr_sdram_s1_end_xfer,
      ddr_sdram_s1_address => ddr_sdram_s1_address,
      ddr_sdram_s1_beginbursttransfer => ddr_sdram_s1_beginbursttransfer,
      ddr_sdram_s1_burstcount => ddr_sdram_s1_burstcount,
      ddr_sdram_s1_byteenable => ddr_sdram_s1_byteenable,
      ddr_sdram_s1_read => ddr_sdram_s1_read,
      ddr_sdram_s1_readdata_from_sa => ddr_sdram_s1_readdata_from_sa,
      ddr_sdram_s1_resetrequest_n_from_sa => ddr_sdram_s1_resetrequest_n_from_sa,
      ddr_sdram_s1_waitrequest_n_from_sa => ddr_sdram_s1_waitrequest_n_from_sa,
      ddr_sdram_s1_write => ddr_sdram_s1_write,
      ddr_sdram_s1_writedata => ddr_sdram_s1_writedata,
      clk => internal_ddr_sdram_phy_clk_out,
      cpu_ddr_clock_bridge_m1_address_to_slave => cpu_ddr_clock_bridge_m1_address_to_slave,
      cpu_ddr_clock_bridge_m1_byteenable => cpu_ddr_clock_bridge_m1_byteenable,
      cpu_ddr_clock_bridge_m1_latency_counter => cpu_ddr_clock_bridge_m1_latency_counter,
      cpu_ddr_clock_bridge_m1_read => cpu_ddr_clock_bridge_m1_read,
      cpu_ddr_clock_bridge_m1_write => cpu_ddr_clock_bridge_m1_write,
      cpu_ddr_clock_bridge_m1_writedata => cpu_ddr_clock_bridge_m1_writedata,
      ddr_sdram_s1_readdata => ddr_sdram_s1_readdata,
      ddr_sdram_s1_readdatavalid => ddr_sdram_s1_readdatavalid,
      ddr_sdram_s1_resetrequest_n => ddr_sdram_s1_resetrequest_n,
      ddr_sdram_s1_waitrequest_n => ddr_sdram_s1_waitrequest_n,
      reset_n => ddr_sdram_phy_clk_out_reset_n
    );


  --ddr_sdram_aux_full_rate_clk_out out_clk assignment, which is an e_assign
  ddr_sdram_aux_full_rate_clk_out <= out_clk_ddr_sdram_aux_full_rate_clk;
  --ddr_sdram_aux_half_rate_clk_out out_clk assignment, which is an e_assign
  ddr_sdram_aux_half_rate_clk_out <= out_clk_ddr_sdram_aux_half_rate_clk;
  --ddr_sdram_phy_clk_out out_clk assignment, which is an e_assign
  internal_ddr_sdram_phy_clk_out <= out_clk_ddr_sdram_phy_clk;
  --reset is asserted asynchronously and deasserted synchronously
  gpib_edm1_reset_clk_0_domain_synch : gpib_edm1_reset_clk_0_domain_synch_module
    port map(
      data_out => clk_0_reset_n,
      clk => clk_0,
      data_in => module_input15,
      reset_n => reset_n_sources
    );

  module_input15 <= std_logic'('1');

  --reset sources mux, which is an e_mux
  reset_n_sources <= Vector_To_Std_Logic(NOT (((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT reset_n))) OR std_logic_vector'("00000000000000000000000000000000")) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_0_jtag_debug_module_resetrequest_from_sa)))) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT ddr_sdram_s1_resetrequest_n_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT ddr_sdram_s1_resetrequest_n_from_sa)))) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pll_s1_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pll_s1_resetrequest_from_sa)))) OR std_logic_vector'("00000000000000000000000000000000"))));
  --the_ddr_sdram, which is an e_ptf_instance
  the_ddr_sdram : ddr_sdram
    port map(
      aux_full_rate_clk => out_clk_ddr_sdram_aux_full_rate_clk,
      aux_half_rate_clk => out_clk_ddr_sdram_aux_half_rate_clk,
      local_init_done => internal_local_init_done_from_the_ddr_sdram,
      local_rdata => ddr_sdram_s1_readdata,
      local_rdata_valid => ddr_sdram_s1_readdatavalid,
      local_ready => ddr_sdram_s1_waitrequest_n,
      local_refresh_ack => internal_local_refresh_ack_from_the_ddr_sdram,
      local_wdata_req => internal_local_wdata_req_from_the_ddr_sdram,
      mem_addr => internal_mem_addr_from_the_ddr_sdram,
      mem_ba => internal_mem_ba_from_the_ddr_sdram,
      mem_cas_n => internal_mem_cas_n_from_the_ddr_sdram,
      mem_cke(0) => internal_mem_cke_from_the_ddr_sdram,
      mem_clk(0) => mem_clk_to_and_from_the_ddr_sdram,
      mem_clk_n(0) => mem_clk_n_to_and_from_the_ddr_sdram,
      mem_cs_n(0) => internal_mem_cs_n_from_the_ddr_sdram,
      mem_dm => internal_mem_dm_from_the_ddr_sdram,
      mem_dq => mem_dq_to_and_from_the_ddr_sdram,
      mem_dqs => mem_dqs_to_and_from_the_ddr_sdram,
      mem_ras_n => internal_mem_ras_n_from_the_ddr_sdram,
      mem_we_n => internal_mem_we_n_from_the_ddr_sdram,
      phy_clk => out_clk_ddr_sdram_phy_clk,
      reset_phy_clk_n => internal_reset_phy_clk_n_from_the_ddr_sdram,
      reset_request_n => ddr_sdram_s1_resetrequest_n,
      global_reset_n => global_reset_n_to_the_ddr_sdram,
      local_address => ddr_sdram_s1_address,
      local_be => ddr_sdram_s1_byteenable,
      local_burstbegin => ddr_sdram_s1_beginbursttransfer,
      local_read_req => ddr_sdram_s1_read,
      local_size => ddr_sdram_s1_burstcount,
      local_wdata => ddr_sdram_s1_writedata,
      local_write_req => ddr_sdram_s1_write,
      pll_ref_clk => clk_0,
      soft_reset_n => clk_0_reset_n
    );


  --the_flash_ssram_pipeline_bridge_s1, which is an e_instance
  the_flash_ssram_pipeline_bridge_s1 : flash_ssram_pipeline_bridge_s1_arbitrator
    port map(
      cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1 => cpu_0_data_master_granted_flash_ssram_pipeline_bridge_s1,
      cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1 => cpu_0_data_master_qualified_request_flash_ssram_pipeline_bridge_s1,
      cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1 => cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1,
      cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register => cpu_0_data_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
      cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1 => cpu_0_data_master_requests_flash_ssram_pipeline_bridge_s1,
      cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1 => cpu_0_instruction_master_granted_flash_ssram_pipeline_bridge_s1,
      cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1 => cpu_0_instruction_master_qualified_request_flash_ssram_pipeline_bridge_s1,
      cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1 => cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1,
      cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register => cpu_0_instruction_master_read_data_valid_flash_ssram_pipeline_bridge_s1_shift_register,
      cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1 => cpu_0_instruction_master_requests_flash_ssram_pipeline_bridge_s1,
      d1_flash_ssram_pipeline_bridge_s1_end_xfer => d1_flash_ssram_pipeline_bridge_s1_end_xfer,
      flash_ssram_pipeline_bridge_s1_address => flash_ssram_pipeline_bridge_s1_address,
      flash_ssram_pipeline_bridge_s1_arbiterlock => flash_ssram_pipeline_bridge_s1_arbiterlock,
      flash_ssram_pipeline_bridge_s1_arbiterlock2 => flash_ssram_pipeline_bridge_s1_arbiterlock2,
      flash_ssram_pipeline_bridge_s1_burstcount => flash_ssram_pipeline_bridge_s1_burstcount,
      flash_ssram_pipeline_bridge_s1_byteenable => flash_ssram_pipeline_bridge_s1_byteenable,
      flash_ssram_pipeline_bridge_s1_chipselect => flash_ssram_pipeline_bridge_s1_chipselect,
      flash_ssram_pipeline_bridge_s1_debugaccess => flash_ssram_pipeline_bridge_s1_debugaccess,
      flash_ssram_pipeline_bridge_s1_endofpacket_from_sa => flash_ssram_pipeline_bridge_s1_endofpacket_from_sa,
      flash_ssram_pipeline_bridge_s1_nativeaddress => flash_ssram_pipeline_bridge_s1_nativeaddress,
      flash_ssram_pipeline_bridge_s1_read => flash_ssram_pipeline_bridge_s1_read,
      flash_ssram_pipeline_bridge_s1_readdata_from_sa => flash_ssram_pipeline_bridge_s1_readdata_from_sa,
      flash_ssram_pipeline_bridge_s1_reset_n => flash_ssram_pipeline_bridge_s1_reset_n,
      flash_ssram_pipeline_bridge_s1_waitrequest_from_sa => flash_ssram_pipeline_bridge_s1_waitrequest_from_sa,
      flash_ssram_pipeline_bridge_s1_write => flash_ssram_pipeline_bridge_s1_write,
      flash_ssram_pipeline_bridge_s1_writedata => flash_ssram_pipeline_bridge_s1_writedata,
      clk => internal_cpu_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_debugaccess => cpu_0_data_master_debugaccess,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_waitrequest => cpu_0_data_master_waitrequest,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      cpu_0_instruction_master_address_to_slave => cpu_0_instruction_master_address_to_slave,
      cpu_0_instruction_master_read => cpu_0_instruction_master_read,
      flash_ssram_pipeline_bridge_s1_endofpacket => flash_ssram_pipeline_bridge_s1_endofpacket,
      flash_ssram_pipeline_bridge_s1_readdata => flash_ssram_pipeline_bridge_s1_readdata,
      flash_ssram_pipeline_bridge_s1_readdatavalid => flash_ssram_pipeline_bridge_s1_readdatavalid,
      flash_ssram_pipeline_bridge_s1_waitrequest => flash_ssram_pipeline_bridge_s1_waitrequest,
      reset_n => cpu_clk_reset_n
    );


  --the_flash_ssram_pipeline_bridge_m1, which is an e_instance
  the_flash_ssram_pipeline_bridge_m1 : flash_ssram_pipeline_bridge_m1_arbitrator
    port map(
      flash_ssram_pipeline_bridge_m1_address_to_slave => flash_ssram_pipeline_bridge_m1_address_to_slave,
      flash_ssram_pipeline_bridge_m1_endofpacket => flash_ssram_pipeline_bridge_m1_endofpacket,
      flash_ssram_pipeline_bridge_m1_latency_counter => flash_ssram_pipeline_bridge_m1_latency_counter,
      flash_ssram_pipeline_bridge_m1_readdata => flash_ssram_pipeline_bridge_m1_readdata,
      flash_ssram_pipeline_bridge_m1_readdatavalid => flash_ssram_pipeline_bridge_m1_readdatavalid,
      flash_ssram_pipeline_bridge_m1_waitrequest => flash_ssram_pipeline_bridge_m1_waitrequest,
      clk => internal_cpu_clk,
      d1_pipeline_bridge_before_tristate_s1_end_xfer => d1_pipeline_bridge_before_tristate_s1_end_xfer,
      flash_ssram_pipeline_bridge_m1_address => flash_ssram_pipeline_bridge_m1_address,
      flash_ssram_pipeline_bridge_m1_burstcount => flash_ssram_pipeline_bridge_m1_burstcount,
      flash_ssram_pipeline_bridge_m1_byteenable => flash_ssram_pipeline_bridge_m1_byteenable,
      flash_ssram_pipeline_bridge_m1_chipselect => flash_ssram_pipeline_bridge_m1_chipselect,
      flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 => flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1,
      flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 => flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1,
      flash_ssram_pipeline_bridge_m1_read => flash_ssram_pipeline_bridge_m1_read,
      flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1 => flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1,
      flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1_shift_register => flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1_shift_register,
      flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 => flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1,
      flash_ssram_pipeline_bridge_m1_write => flash_ssram_pipeline_bridge_m1_write,
      flash_ssram_pipeline_bridge_m1_writedata => flash_ssram_pipeline_bridge_m1_writedata,
      pipeline_bridge_before_tristate_s1_endofpacket_from_sa => pipeline_bridge_before_tristate_s1_endofpacket_from_sa,
      pipeline_bridge_before_tristate_s1_readdata_from_sa => pipeline_bridge_before_tristate_s1_readdata_from_sa,
      pipeline_bridge_before_tristate_s1_waitrequest_from_sa => pipeline_bridge_before_tristate_s1_waitrequest_from_sa,
      reset_n => cpu_clk_reset_n
    );


  --the_flash_ssram_pipeline_bridge, which is an e_ptf_instance
  the_flash_ssram_pipeline_bridge : flash_ssram_pipeline_bridge
    port map(
      m1_address => flash_ssram_pipeline_bridge_m1_address,
      m1_burstcount => flash_ssram_pipeline_bridge_m1_burstcount,
      m1_byteenable => flash_ssram_pipeline_bridge_m1_byteenable,
      m1_chipselect => flash_ssram_pipeline_bridge_m1_chipselect,
      m1_debugaccess => flash_ssram_pipeline_bridge_m1_debugaccess,
      m1_read => flash_ssram_pipeline_bridge_m1_read,
      m1_write => flash_ssram_pipeline_bridge_m1_write,
      m1_writedata => flash_ssram_pipeline_bridge_m1_writedata,
      s1_endofpacket => flash_ssram_pipeline_bridge_s1_endofpacket,
      s1_readdata => flash_ssram_pipeline_bridge_s1_readdata,
      s1_readdatavalid => flash_ssram_pipeline_bridge_s1_readdatavalid,
      s1_waitrequest => flash_ssram_pipeline_bridge_s1_waitrequest,
      clk => internal_cpu_clk,
      m1_endofpacket => flash_ssram_pipeline_bridge_m1_endofpacket,
      m1_readdata => flash_ssram_pipeline_bridge_m1_readdata,
      m1_readdatavalid => flash_ssram_pipeline_bridge_m1_readdatavalid,
      m1_waitrequest => flash_ssram_pipeline_bridge_m1_waitrequest,
      reset_n => flash_ssram_pipeline_bridge_s1_reset_n,
      s1_address => flash_ssram_pipeline_bridge_s1_address,
      s1_arbiterlock => flash_ssram_pipeline_bridge_s1_arbiterlock,
      s1_arbiterlock2 => flash_ssram_pipeline_bridge_s1_arbiterlock2,
      s1_burstcount => flash_ssram_pipeline_bridge_s1_burstcount,
      s1_byteenable => flash_ssram_pipeline_bridge_s1_byteenable,
      s1_chipselect => flash_ssram_pipeline_bridge_s1_chipselect,
      s1_debugaccess => flash_ssram_pipeline_bridge_s1_debugaccess,
      s1_nativeaddress => flash_ssram_pipeline_bridge_s1_nativeaddress,
      s1_read => flash_ssram_pipeline_bridge_s1_read,
      s1_write => flash_ssram_pipeline_bridge_s1_write,
      s1_writedata => flash_ssram_pipeline_bridge_s1_writedata
    );


  --the_flash_ssram_tristate_avalon_slave, which is an e_instance
  the_flash_ssram_tristate_avalon_slave : flash_ssram_tristate_avalon_slave_arbitrator
    port map(
      adsc_n_to_the_ssram => internal_adsc_n_to_the_ssram,
      bw_n_to_the_ssram => internal_bw_n_to_the_ssram,
      bwe_n_to_the_ssram => internal_bwe_n_to_the_ssram,
      cfi_flash_s1_wait_counter_eq_0 => cfi_flash_s1_wait_counter_eq_0,
      chipenable1_n_to_the_ssram => internal_chipenable1_n_to_the_ssram,
      d1_flash_ssram_tristate_avalon_slave_end_xfer => d1_flash_ssram_tristate_avalon_slave_end_xfer,
      flash_ssram_tristate_address => internal_flash_ssram_tristate_address,
      flash_ssram_tristate_data => flash_ssram_tristate_data,
      incoming_flash_ssram_tristate_data => incoming_flash_ssram_tristate_data,
      incoming_flash_ssram_tristate_data_with_Xs_converted_to_0 => incoming_flash_ssram_tristate_data_with_Xs_converted_to_0,
      outputenable_n_to_the_ssram => internal_outputenable_n_to_the_ssram,
      pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1 => pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1,
      pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 => pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1,
      pipeline_bridge_before_tristate_m1_granted_ssram_s1 => pipeline_bridge_before_tristate_m1_granted_ssram_s1,
      pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 => pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1,
      pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 => pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1,
      pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1 => pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1,
      pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1 => pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1,
      pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 => pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1,
      pipeline_bridge_before_tristate_m1_requests_ssram_s1 => pipeline_bridge_before_tristate_m1_requests_ssram_s1,
      read_n_to_the_cfi_flash => internal_read_n_to_the_cfi_flash,
      reset_n_to_the_ssram => internal_reset_n_to_the_ssram,
      select_n_to_the_cfi_flash => internal_select_n_to_the_cfi_flash,
      write_n_to_the_cfi_flash => internal_write_n_to_the_cfi_flash,
      clk => internal_cpu_clk,
      pipeline_bridge_before_tristate_m1_address_to_slave => pipeline_bridge_before_tristate_m1_address_to_slave,
      pipeline_bridge_before_tristate_m1_burstcount => pipeline_bridge_before_tristate_m1_burstcount,
      pipeline_bridge_before_tristate_m1_byteenable => pipeline_bridge_before_tristate_m1_byteenable,
      pipeline_bridge_before_tristate_m1_chipselect => pipeline_bridge_before_tristate_m1_chipselect,
      pipeline_bridge_before_tristate_m1_dbs_address => pipeline_bridge_before_tristate_m1_dbs_address,
      pipeline_bridge_before_tristate_m1_dbs_write_16 => pipeline_bridge_before_tristate_m1_dbs_write_16,
      pipeline_bridge_before_tristate_m1_latency_counter => pipeline_bridge_before_tristate_m1_latency_counter,
      pipeline_bridge_before_tristate_m1_read => pipeline_bridge_before_tristate_m1_read,
      pipeline_bridge_before_tristate_m1_write => pipeline_bridge_before_tristate_m1_write,
      pipeline_bridge_before_tristate_m1_writedata => pipeline_bridge_before_tristate_m1_writedata,
      reset_n => cpu_clk_reset_n
    );


  --the_gpib_edm1_clock_0_in, which is an e_instance
  the_gpib_edm1_clock_0_in : gpib_edm1_clock_0_in_arbitrator
    port map(
      cpu_0_data_master_granted_gpib_edm1_clock_0_in => cpu_0_data_master_granted_gpib_edm1_clock_0_in,
      cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in => cpu_0_data_master_qualified_request_gpib_edm1_clock_0_in,
      cpu_0_data_master_read_data_valid_gpib_edm1_clock_0_in => cpu_0_data_master_read_data_valid_gpib_edm1_clock_0_in,
      cpu_0_data_master_requests_gpib_edm1_clock_0_in => cpu_0_data_master_requests_gpib_edm1_clock_0_in,
      d1_gpib_edm1_clock_0_in_end_xfer => d1_gpib_edm1_clock_0_in_end_xfer,
      gpib_edm1_clock_0_in_address => gpib_edm1_clock_0_in_address,
      gpib_edm1_clock_0_in_byteenable => gpib_edm1_clock_0_in_byteenable,
      gpib_edm1_clock_0_in_endofpacket_from_sa => gpib_edm1_clock_0_in_endofpacket_from_sa,
      gpib_edm1_clock_0_in_nativeaddress => gpib_edm1_clock_0_in_nativeaddress,
      gpib_edm1_clock_0_in_read => gpib_edm1_clock_0_in_read,
      gpib_edm1_clock_0_in_readdata_from_sa => gpib_edm1_clock_0_in_readdata_from_sa,
      gpib_edm1_clock_0_in_reset_n => gpib_edm1_clock_0_in_reset_n,
      gpib_edm1_clock_0_in_waitrequest_from_sa => gpib_edm1_clock_0_in_waitrequest_from_sa,
      gpib_edm1_clock_0_in_write => gpib_edm1_clock_0_in_write,
      gpib_edm1_clock_0_in_writedata => gpib_edm1_clock_0_in_writedata,
      clk => internal_cpu_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_waitrequest => cpu_0_data_master_waitrequest,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      gpib_edm1_clock_0_in_endofpacket => gpib_edm1_clock_0_in_endofpacket,
      gpib_edm1_clock_0_in_readdata => gpib_edm1_clock_0_in_readdata,
      gpib_edm1_clock_0_in_waitrequest => gpib_edm1_clock_0_in_waitrequest,
      reset_n => cpu_clk_reset_n
    );


  --the_gpib_edm1_clock_0_out, which is an e_instance
  the_gpib_edm1_clock_0_out : gpib_edm1_clock_0_out_arbitrator
    port map(
      gpib_edm1_clock_0_out_address_to_slave => gpib_edm1_clock_0_out_address_to_slave,
      gpib_edm1_clock_0_out_readdata => gpib_edm1_clock_0_out_readdata,
      gpib_edm1_clock_0_out_reset_n => gpib_edm1_clock_0_out_reset_n,
      gpib_edm1_clock_0_out_waitrequest => gpib_edm1_clock_0_out_waitrequest,
      clk => clk_0,
      d1_pll_s1_end_xfer => d1_pll_s1_end_xfer,
      gpib_edm1_clock_0_out_address => gpib_edm1_clock_0_out_address,
      gpib_edm1_clock_0_out_byteenable => gpib_edm1_clock_0_out_byteenable,
      gpib_edm1_clock_0_out_granted_pll_s1 => gpib_edm1_clock_0_out_granted_pll_s1,
      gpib_edm1_clock_0_out_qualified_request_pll_s1 => gpib_edm1_clock_0_out_qualified_request_pll_s1,
      gpib_edm1_clock_0_out_read => gpib_edm1_clock_0_out_read,
      gpib_edm1_clock_0_out_read_data_valid_pll_s1 => gpib_edm1_clock_0_out_read_data_valid_pll_s1,
      gpib_edm1_clock_0_out_requests_pll_s1 => gpib_edm1_clock_0_out_requests_pll_s1,
      gpib_edm1_clock_0_out_write => gpib_edm1_clock_0_out_write,
      gpib_edm1_clock_0_out_writedata => gpib_edm1_clock_0_out_writedata,
      pll_s1_readdata_from_sa => pll_s1_readdata_from_sa,
      reset_n => clk_0_reset_n
    );


  --the_gpib_edm1_clock_0, which is an e_ptf_instance
  the_gpib_edm1_clock_0 : gpib_edm1_clock_0
    port map(
      master_address => gpib_edm1_clock_0_out_address,
      master_byteenable => gpib_edm1_clock_0_out_byteenable,
      master_nativeaddress => gpib_edm1_clock_0_out_nativeaddress,
      master_read => gpib_edm1_clock_0_out_read,
      master_write => gpib_edm1_clock_0_out_write,
      master_writedata => gpib_edm1_clock_0_out_writedata,
      slave_endofpacket => gpib_edm1_clock_0_in_endofpacket,
      slave_readdata => gpib_edm1_clock_0_in_readdata,
      slave_waitrequest => gpib_edm1_clock_0_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => gpib_edm1_clock_0_out_endofpacket,
      master_readdata => gpib_edm1_clock_0_out_readdata,
      master_reset_n => gpib_edm1_clock_0_out_reset_n,
      master_waitrequest => gpib_edm1_clock_0_out_waitrequest,
      slave_address => gpib_edm1_clock_0_in_address,
      slave_byteenable => gpib_edm1_clock_0_in_byteenable,
      slave_clk => internal_cpu_clk,
      slave_nativeaddress => gpib_edm1_clock_0_in_nativeaddress,
      slave_read => gpib_edm1_clock_0_in_read,
      slave_reset_n => gpib_edm1_clock_0_in_reset_n,
      slave_write => gpib_edm1_clock_0_in_write,
      slave_writedata => gpib_edm1_clock_0_in_writedata
    );


  --the_gpib_edm1_clock_1_in, which is an e_instance
  the_gpib_edm1_clock_1_in : gpib_edm1_clock_1_in_arbitrator
    port map(
      cpu_0_data_master_granted_gpib_edm1_clock_1_in => cpu_0_data_master_granted_gpib_edm1_clock_1_in,
      cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in => cpu_0_data_master_qualified_request_gpib_edm1_clock_1_in,
      cpu_0_data_master_read_data_valid_gpib_edm1_clock_1_in => cpu_0_data_master_read_data_valid_gpib_edm1_clock_1_in,
      cpu_0_data_master_requests_gpib_edm1_clock_1_in => cpu_0_data_master_requests_gpib_edm1_clock_1_in,
      d1_gpib_edm1_clock_1_in_end_xfer => d1_gpib_edm1_clock_1_in_end_xfer,
      gpib_edm1_clock_1_in_address => gpib_edm1_clock_1_in_address,
      gpib_edm1_clock_1_in_byteenable => gpib_edm1_clock_1_in_byteenable,
      gpib_edm1_clock_1_in_endofpacket_from_sa => gpib_edm1_clock_1_in_endofpacket_from_sa,
      gpib_edm1_clock_1_in_nativeaddress => gpib_edm1_clock_1_in_nativeaddress,
      gpib_edm1_clock_1_in_read => gpib_edm1_clock_1_in_read,
      gpib_edm1_clock_1_in_readdata_from_sa => gpib_edm1_clock_1_in_readdata_from_sa,
      gpib_edm1_clock_1_in_reset_n => gpib_edm1_clock_1_in_reset_n,
      gpib_edm1_clock_1_in_waitrequest_from_sa => gpib_edm1_clock_1_in_waitrequest_from_sa,
      gpib_edm1_clock_1_in_write => gpib_edm1_clock_1_in_write,
      gpib_edm1_clock_1_in_writedata => gpib_edm1_clock_1_in_writedata,
      clk => internal_cpu_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_waitrequest => cpu_0_data_master_waitrequest,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      gpib_edm1_clock_1_in_endofpacket => gpib_edm1_clock_1_in_endofpacket,
      gpib_edm1_clock_1_in_readdata => gpib_edm1_clock_1_in_readdata,
      gpib_edm1_clock_1_in_waitrequest => gpib_edm1_clock_1_in_waitrequest,
      reset_n => cpu_clk_reset_n
    );


  --the_gpib_edm1_clock_1_out, which is an e_instance
  the_gpib_edm1_clock_1_out : gpib_edm1_clock_1_out_arbitrator
    port map(
      gpib_edm1_clock_1_out_address_to_slave => gpib_edm1_clock_1_out_address_to_slave,
      gpib_edm1_clock_1_out_readdata => gpib_edm1_clock_1_out_readdata,
      gpib_edm1_clock_1_out_reset_n => gpib_edm1_clock_1_out_reset_n,
      gpib_edm1_clock_1_out_waitrequest => gpib_edm1_clock_1_out_waitrequest,
      clk => internal_pll_c3_out,
      d1_remote_update_cycloneiii_1_s1_end_xfer => d1_remote_update_cycloneiii_1_s1_end_xfer,
      gpib_edm1_clock_1_out_address => gpib_edm1_clock_1_out_address,
      gpib_edm1_clock_1_out_byteenable => gpib_edm1_clock_1_out_byteenable,
      gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 => gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1,
      gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 => gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1,
      gpib_edm1_clock_1_out_read => gpib_edm1_clock_1_out_read,
      gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1 => gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1,
      gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 => gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1,
      gpib_edm1_clock_1_out_write => gpib_edm1_clock_1_out_write,
      gpib_edm1_clock_1_out_writedata => gpib_edm1_clock_1_out_writedata,
      remote_update_cycloneiii_1_s1_readdata_from_sa => remote_update_cycloneiii_1_s1_readdata_from_sa,
      remote_update_cycloneiii_1_s1_waitrequest_from_sa => remote_update_cycloneiii_1_s1_waitrequest_from_sa,
      reset_n => pll_c3_out_reset_n
    );


  --the_gpib_edm1_clock_1, which is an e_ptf_instance
  the_gpib_edm1_clock_1 : gpib_edm1_clock_1
    port map(
      master_address => gpib_edm1_clock_1_out_address,
      master_byteenable => gpib_edm1_clock_1_out_byteenable,
      master_nativeaddress => gpib_edm1_clock_1_out_nativeaddress,
      master_read => gpib_edm1_clock_1_out_read,
      master_write => gpib_edm1_clock_1_out_write,
      master_writedata => gpib_edm1_clock_1_out_writedata,
      slave_endofpacket => gpib_edm1_clock_1_in_endofpacket,
      slave_readdata => gpib_edm1_clock_1_in_readdata,
      slave_waitrequest => gpib_edm1_clock_1_in_waitrequest,
      master_clk => internal_pll_c3_out,
      master_endofpacket => gpib_edm1_clock_1_out_endofpacket,
      master_readdata => gpib_edm1_clock_1_out_readdata,
      master_reset_n => gpib_edm1_clock_1_out_reset_n,
      master_waitrequest => gpib_edm1_clock_1_out_waitrequest,
      slave_address => gpib_edm1_clock_1_in_address,
      slave_byteenable => gpib_edm1_clock_1_in_byteenable,
      slave_clk => internal_cpu_clk,
      slave_nativeaddress => gpib_edm1_clock_1_in_nativeaddress,
      slave_read => gpib_edm1_clock_1_in_read,
      slave_reset_n => gpib_edm1_clock_1_in_reset_n,
      slave_write => gpib_edm1_clock_1_in_write,
      slave_writedata => gpib_edm1_clock_1_in_writedata
    );


  --the_gpib_edm1_clock_2_in, which is an e_instance
  the_gpib_edm1_clock_2_in : gpib_edm1_clock_2_in_arbitrator
    port map(
      clock_crossing_0_m1_granted_gpib_edm1_clock_2_in => clock_crossing_0_m1_granted_gpib_edm1_clock_2_in,
      clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in => clock_crossing_0_m1_qualified_request_gpib_edm1_clock_2_in,
      clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in => clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_2_in,
      clock_crossing_0_m1_requests_gpib_edm1_clock_2_in => clock_crossing_0_m1_requests_gpib_edm1_clock_2_in,
      d1_gpib_edm1_clock_2_in_end_xfer => d1_gpib_edm1_clock_2_in_end_xfer,
      gpib_edm1_clock_2_in_address => gpib_edm1_clock_2_in_address,
      gpib_edm1_clock_2_in_byteenable => gpib_edm1_clock_2_in_byteenable,
      gpib_edm1_clock_2_in_endofpacket_from_sa => gpib_edm1_clock_2_in_endofpacket_from_sa,
      gpib_edm1_clock_2_in_nativeaddress => gpib_edm1_clock_2_in_nativeaddress,
      gpib_edm1_clock_2_in_read => gpib_edm1_clock_2_in_read,
      gpib_edm1_clock_2_in_readdata_from_sa => gpib_edm1_clock_2_in_readdata_from_sa,
      gpib_edm1_clock_2_in_reset_n => gpib_edm1_clock_2_in_reset_n,
      gpib_edm1_clock_2_in_waitrequest_from_sa => gpib_edm1_clock_2_in_waitrequest_from_sa,
      gpib_edm1_clock_2_in_write => gpib_edm1_clock_2_in_write,
      gpib_edm1_clock_2_in_writedata => gpib_edm1_clock_2_in_writedata,
      clk => internal_pll_c2_out,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_byteenable => clock_crossing_0_m1_byteenable,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      gpib_edm1_clock_2_in_endofpacket => gpib_edm1_clock_2_in_endofpacket,
      gpib_edm1_clock_2_in_readdata => gpib_edm1_clock_2_in_readdata,
      gpib_edm1_clock_2_in_waitrequest => gpib_edm1_clock_2_in_waitrequest,
      reset_n => pll_c2_out_reset_n
    );


  --the_gpib_edm1_clock_2_out, which is an e_instance
  the_gpib_edm1_clock_2_out : gpib_edm1_clock_2_out_arbitrator
    port map(
      gpib_edm1_clock_2_out_address_to_slave => gpib_edm1_clock_2_out_address_to_slave,
      gpib_edm1_clock_2_out_endofpacket => gpib_edm1_clock_2_out_endofpacket,
      gpib_edm1_clock_2_out_readdata => gpib_edm1_clock_2_out_readdata,
      gpib_edm1_clock_2_out_reset_n => gpib_edm1_clock_2_out_reset_n,
      gpib_edm1_clock_2_out_waitrequest => gpib_edm1_clock_2_out_waitrequest,
      ad7928_spi_control_port_endofpacket_from_sa => ad7928_spi_control_port_endofpacket_from_sa,
      ad7928_spi_control_port_readdata_from_sa => ad7928_spi_control_port_readdata_from_sa,
      clk => internal_cpu_clk,
      d1_ad7928_spi_control_port_end_xfer => d1_ad7928_spi_control_port_end_xfer,
      gpib_edm1_clock_2_out_address => gpib_edm1_clock_2_out_address,
      gpib_edm1_clock_2_out_byteenable => gpib_edm1_clock_2_out_byteenable,
      gpib_edm1_clock_2_out_granted_ad7928_spi_control_port => gpib_edm1_clock_2_out_granted_ad7928_spi_control_port,
      gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port => gpib_edm1_clock_2_out_qualified_request_ad7928_spi_control_port,
      gpib_edm1_clock_2_out_read => gpib_edm1_clock_2_out_read,
      gpib_edm1_clock_2_out_read_data_valid_ad7928_spi_control_port => gpib_edm1_clock_2_out_read_data_valid_ad7928_spi_control_port,
      gpib_edm1_clock_2_out_requests_ad7928_spi_control_port => gpib_edm1_clock_2_out_requests_ad7928_spi_control_port,
      gpib_edm1_clock_2_out_write => gpib_edm1_clock_2_out_write,
      gpib_edm1_clock_2_out_writedata => gpib_edm1_clock_2_out_writedata,
      reset_n => cpu_clk_reset_n
    );


  --the_gpib_edm1_clock_2, which is an e_ptf_instance
  the_gpib_edm1_clock_2 : gpib_edm1_clock_2
    port map(
      master_address => gpib_edm1_clock_2_out_address,
      master_byteenable => gpib_edm1_clock_2_out_byteenable,
      master_nativeaddress => gpib_edm1_clock_2_out_nativeaddress,
      master_read => gpib_edm1_clock_2_out_read,
      master_write => gpib_edm1_clock_2_out_write,
      master_writedata => gpib_edm1_clock_2_out_writedata,
      slave_endofpacket => gpib_edm1_clock_2_in_endofpacket,
      slave_readdata => gpib_edm1_clock_2_in_readdata,
      slave_waitrequest => gpib_edm1_clock_2_in_waitrequest,
      master_clk => internal_cpu_clk,
      master_endofpacket => gpib_edm1_clock_2_out_endofpacket,
      master_readdata => gpib_edm1_clock_2_out_readdata,
      master_reset_n => gpib_edm1_clock_2_out_reset_n,
      master_waitrequest => gpib_edm1_clock_2_out_waitrequest,
      slave_address => gpib_edm1_clock_2_in_address,
      slave_byteenable => gpib_edm1_clock_2_in_byteenable,
      slave_clk => internal_pll_c2_out,
      slave_nativeaddress => gpib_edm1_clock_2_in_nativeaddress,
      slave_read => gpib_edm1_clock_2_in_read,
      slave_reset_n => gpib_edm1_clock_2_in_reset_n,
      slave_write => gpib_edm1_clock_2_in_write,
      slave_writedata => gpib_edm1_clock_2_in_writedata
    );


  --the_gpib_edm1_clock_3_in, which is an e_instance
  the_gpib_edm1_clock_3_in : gpib_edm1_clock_3_in_arbitrator
    port map(
      clock_crossing_0_m1_granted_gpib_edm1_clock_3_in => clock_crossing_0_m1_granted_gpib_edm1_clock_3_in,
      clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in => clock_crossing_0_m1_qualified_request_gpib_edm1_clock_3_in,
      clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in => clock_crossing_0_m1_read_data_valid_gpib_edm1_clock_3_in,
      clock_crossing_0_m1_requests_gpib_edm1_clock_3_in => clock_crossing_0_m1_requests_gpib_edm1_clock_3_in,
      d1_gpib_edm1_clock_3_in_end_xfer => d1_gpib_edm1_clock_3_in_end_xfer,
      gpib_edm1_clock_3_in_address => gpib_edm1_clock_3_in_address,
      gpib_edm1_clock_3_in_byteenable => gpib_edm1_clock_3_in_byteenable,
      gpib_edm1_clock_3_in_endofpacket_from_sa => gpib_edm1_clock_3_in_endofpacket_from_sa,
      gpib_edm1_clock_3_in_nativeaddress => gpib_edm1_clock_3_in_nativeaddress,
      gpib_edm1_clock_3_in_read => gpib_edm1_clock_3_in_read,
      gpib_edm1_clock_3_in_readdata_from_sa => gpib_edm1_clock_3_in_readdata_from_sa,
      gpib_edm1_clock_3_in_reset_n => gpib_edm1_clock_3_in_reset_n,
      gpib_edm1_clock_3_in_waitrequest_from_sa => gpib_edm1_clock_3_in_waitrequest_from_sa,
      gpib_edm1_clock_3_in_write => gpib_edm1_clock_3_in_write,
      gpib_edm1_clock_3_in_writedata => gpib_edm1_clock_3_in_writedata,
      clk => internal_pll_c2_out,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_byteenable => clock_crossing_0_m1_byteenable,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      gpib_edm1_clock_3_in_endofpacket => gpib_edm1_clock_3_in_endofpacket,
      gpib_edm1_clock_3_in_readdata => gpib_edm1_clock_3_in_readdata,
      gpib_edm1_clock_3_in_waitrequest => gpib_edm1_clock_3_in_waitrequest,
      reset_n => pll_c2_out_reset_n
    );


  --the_gpib_edm1_clock_3_out, which is an e_instance
  the_gpib_edm1_clock_3_out : gpib_edm1_clock_3_out_arbitrator
    port map(
      gpib_edm1_clock_3_out_address_to_slave => gpib_edm1_clock_3_out_address_to_slave,
      gpib_edm1_clock_3_out_endofpacket => gpib_edm1_clock_3_out_endofpacket,
      gpib_edm1_clock_3_out_readdata => gpib_edm1_clock_3_out_readdata,
      gpib_edm1_clock_3_out_reset_n => gpib_edm1_clock_3_out_reset_n,
      gpib_edm1_clock_3_out_waitrequest => gpib_edm1_clock_3_out_waitrequest,
      clk => internal_cpu_clk,
      d1_dac_ad5308_spi_control_port_end_xfer => d1_dac_ad5308_spi_control_port_end_xfer,
      dac_ad5308_spi_control_port_endofpacket_from_sa => dac_ad5308_spi_control_port_endofpacket_from_sa,
      dac_ad5308_spi_control_port_readdata_from_sa => dac_ad5308_spi_control_port_readdata_from_sa,
      gpib_edm1_clock_3_out_address => gpib_edm1_clock_3_out_address,
      gpib_edm1_clock_3_out_byteenable => gpib_edm1_clock_3_out_byteenable,
      gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port => gpib_edm1_clock_3_out_granted_dac_ad5308_spi_control_port,
      gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port => gpib_edm1_clock_3_out_qualified_request_dac_ad5308_spi_control_port,
      gpib_edm1_clock_3_out_read => gpib_edm1_clock_3_out_read,
      gpib_edm1_clock_3_out_read_data_valid_dac_ad5308_spi_control_port => gpib_edm1_clock_3_out_read_data_valid_dac_ad5308_spi_control_port,
      gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port => gpib_edm1_clock_3_out_requests_dac_ad5308_spi_control_port,
      gpib_edm1_clock_3_out_write => gpib_edm1_clock_3_out_write,
      gpib_edm1_clock_3_out_writedata => gpib_edm1_clock_3_out_writedata,
      reset_n => cpu_clk_reset_n
    );


  --the_gpib_edm1_clock_3, which is an e_ptf_instance
  the_gpib_edm1_clock_3 : gpib_edm1_clock_3
    port map(
      master_address => gpib_edm1_clock_3_out_address,
      master_byteenable => gpib_edm1_clock_3_out_byteenable,
      master_nativeaddress => gpib_edm1_clock_3_out_nativeaddress,
      master_read => gpib_edm1_clock_3_out_read,
      master_write => gpib_edm1_clock_3_out_write,
      master_writedata => gpib_edm1_clock_3_out_writedata,
      slave_endofpacket => gpib_edm1_clock_3_in_endofpacket,
      slave_readdata => gpib_edm1_clock_3_in_readdata,
      slave_waitrequest => gpib_edm1_clock_3_in_waitrequest,
      master_clk => internal_cpu_clk,
      master_endofpacket => gpib_edm1_clock_3_out_endofpacket,
      master_readdata => gpib_edm1_clock_3_out_readdata,
      master_reset_n => gpib_edm1_clock_3_out_reset_n,
      master_waitrequest => gpib_edm1_clock_3_out_waitrequest,
      slave_address => gpib_edm1_clock_3_in_address,
      slave_byteenable => gpib_edm1_clock_3_in_byteenable,
      slave_clk => internal_pll_c2_out,
      slave_nativeaddress => gpib_edm1_clock_3_in_nativeaddress,
      slave_read => gpib_edm1_clock_3_in_read,
      slave_reset_n => gpib_edm1_clock_3_in_reset_n,
      slave_write => gpib_edm1_clock_3_in_write,
      slave_writedata => gpib_edm1_clock_3_in_writedata
    );


  --the_gpib_leds_s1, which is an e_instance
  the_gpib_leds_s1 : gpib_leds_s1_arbitrator
    port map(
      clock_crossing_0_m1_granted_gpib_leds_s1 => clock_crossing_0_m1_granted_gpib_leds_s1,
      clock_crossing_0_m1_qualified_request_gpib_leds_s1 => clock_crossing_0_m1_qualified_request_gpib_leds_s1,
      clock_crossing_0_m1_read_data_valid_gpib_leds_s1 => clock_crossing_0_m1_read_data_valid_gpib_leds_s1,
      clock_crossing_0_m1_requests_gpib_leds_s1 => clock_crossing_0_m1_requests_gpib_leds_s1,
      d1_gpib_leds_s1_end_xfer => d1_gpib_leds_s1_end_xfer,
      gpib_leds_s1_address => gpib_leds_s1_address,
      gpib_leds_s1_chipselect => gpib_leds_s1_chipselect,
      gpib_leds_s1_readdata_from_sa => gpib_leds_s1_readdata_from_sa,
      gpib_leds_s1_reset_n => gpib_leds_s1_reset_n,
      gpib_leds_s1_write_n => gpib_leds_s1_write_n,
      gpib_leds_s1_writedata => gpib_leds_s1_writedata,
      clk => internal_pll_c2_out,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_byteenable => clock_crossing_0_m1_byteenable,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      gpib_leds_s1_readdata => gpib_leds_s1_readdata,
      reset_n => pll_c2_out_reset_n
    );


  --the_gpib_leds, which is an e_ptf_instance
  the_gpib_leds : gpib_leds
    port map(
      out_port => internal_out_port_from_the_gpib_leds,
      readdata => gpib_leds_s1_readdata,
      address => gpib_leds_s1_address,
      chipselect => gpib_leds_s1_chipselect,
      clk => internal_pll_c2_out,
      reset_n => gpib_leds_s1_reset_n,
      write_n => gpib_leds_s1_write_n,
      writedata => gpib_leds_s1_writedata
    );


  --the_gpio1_s1, which is an e_instance
  the_gpio1_s1 : gpio1_s1_arbitrator
    port map(
      clock_crossing_0_m1_granted_gpio1_s1 => clock_crossing_0_m1_granted_gpio1_s1,
      clock_crossing_0_m1_qualified_request_gpio1_s1 => clock_crossing_0_m1_qualified_request_gpio1_s1,
      clock_crossing_0_m1_read_data_valid_gpio1_s1 => clock_crossing_0_m1_read_data_valid_gpio1_s1,
      clock_crossing_0_m1_requests_gpio1_s1 => clock_crossing_0_m1_requests_gpio1_s1,
      d1_gpio1_s1_end_xfer => d1_gpio1_s1_end_xfer,
      gpio1_s1_address => gpio1_s1_address,
      gpio1_s1_chipselect => gpio1_s1_chipselect,
      gpio1_s1_readdata_from_sa => gpio1_s1_readdata_from_sa,
      gpio1_s1_reset_n => gpio1_s1_reset_n,
      gpio1_s1_write_n => gpio1_s1_write_n,
      gpio1_s1_writedata => gpio1_s1_writedata,
      clk => internal_pll_c2_out,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_byteenable => clock_crossing_0_m1_byteenable,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      gpio1_s1_readdata => gpio1_s1_readdata,
      reset_n => pll_c2_out_reset_n
    );


  --the_gpio1, which is an e_ptf_instance
  the_gpio1 : gpio1
    port map(
      bidir_port => bidir_port_to_and_from_the_gpio1,
      readdata => gpio1_s1_readdata,
      address => gpio1_s1_address,
      chipselect => gpio1_s1_chipselect,
      clk => internal_pll_c2_out,
      reset_n => gpio1_s1_reset_n,
      write_n => gpio1_s1_write_n,
      writedata => gpio1_s1_writedata
    );


  --the_gpio2_s1, which is an e_instance
  the_gpio2_s1 : gpio2_s1_arbitrator
    port map(
      clock_crossing_0_m1_granted_gpio2_s1 => clock_crossing_0_m1_granted_gpio2_s1,
      clock_crossing_0_m1_qualified_request_gpio2_s1 => clock_crossing_0_m1_qualified_request_gpio2_s1,
      clock_crossing_0_m1_read_data_valid_gpio2_s1 => clock_crossing_0_m1_read_data_valid_gpio2_s1,
      clock_crossing_0_m1_requests_gpio2_s1 => clock_crossing_0_m1_requests_gpio2_s1,
      d1_gpio2_s1_end_xfer => d1_gpio2_s1_end_xfer,
      gpio2_s1_address => gpio2_s1_address,
      gpio2_s1_chipselect => gpio2_s1_chipselect,
      gpio2_s1_readdata_from_sa => gpio2_s1_readdata_from_sa,
      gpio2_s1_reset_n => gpio2_s1_reset_n,
      gpio2_s1_write_n => gpio2_s1_write_n,
      gpio2_s1_writedata => gpio2_s1_writedata,
      clk => internal_pll_c2_out,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_byteenable => clock_crossing_0_m1_byteenable,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      gpio2_s1_readdata => gpio2_s1_readdata,
      reset_n => pll_c2_out_reset_n
    );


  --the_gpio2, which is an e_ptf_instance
  the_gpio2 : gpio2
    port map(
      out_port => internal_out_port_from_the_gpio2,
      readdata => gpio2_s1_readdata,
      address => gpio2_s1_address,
      chipselect => gpio2_s1_chipselect,
      clk => internal_pll_c2_out,
      reset_n => gpio2_s1_reset_n,
      write_n => gpio2_s1_write_n,
      writedata => gpio2_s1_writedata
    );


  --the_high_res_timer_s1, which is an e_instance
  the_high_res_timer_s1 : high_res_timer_s1_arbitrator
    port map(
      clock_crossing_0_m1_granted_high_res_timer_s1 => clock_crossing_0_m1_granted_high_res_timer_s1,
      clock_crossing_0_m1_qualified_request_high_res_timer_s1 => clock_crossing_0_m1_qualified_request_high_res_timer_s1,
      clock_crossing_0_m1_read_data_valid_high_res_timer_s1 => clock_crossing_0_m1_read_data_valid_high_res_timer_s1,
      clock_crossing_0_m1_requests_high_res_timer_s1 => clock_crossing_0_m1_requests_high_res_timer_s1,
      d1_high_res_timer_s1_end_xfer => d1_high_res_timer_s1_end_xfer,
      high_res_timer_s1_address => high_res_timer_s1_address,
      high_res_timer_s1_chipselect => high_res_timer_s1_chipselect,
      high_res_timer_s1_irq_from_sa => high_res_timer_s1_irq_from_sa,
      high_res_timer_s1_readdata_from_sa => high_res_timer_s1_readdata_from_sa,
      high_res_timer_s1_reset_n => high_res_timer_s1_reset_n,
      high_res_timer_s1_write_n => high_res_timer_s1_write_n,
      high_res_timer_s1_writedata => high_res_timer_s1_writedata,
      clk => internal_pll_c2_out,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      high_res_timer_s1_irq => high_res_timer_s1_irq,
      high_res_timer_s1_readdata => high_res_timer_s1_readdata,
      reset_n => pll_c2_out_reset_n
    );


  --the_high_res_timer, which is an e_ptf_instance
  the_high_res_timer : high_res_timer
    port map(
      irq => high_res_timer_s1_irq,
      readdata => high_res_timer_s1_readdata,
      address => high_res_timer_s1_address,
      chipselect => high_res_timer_s1_chipselect,
      clk => internal_pll_c2_out,
      reset_n => high_res_timer_s1_reset_n,
      write_n => high_res_timer_s1_write_n,
      writedata => high_res_timer_s1_writedata
    );


  --the_jtag_uart_avalon_jtag_slave, which is an e_instance
  the_jtag_uart_avalon_jtag_slave : jtag_uart_avalon_jtag_slave_arbitrator
    port map(
      clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave => clock_crossing_0_m1_granted_jtag_uart_avalon_jtag_slave,
      clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave => clock_crossing_0_m1_qualified_request_jtag_uart_avalon_jtag_slave,
      clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave => clock_crossing_0_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
      clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave => clock_crossing_0_m1_requests_jtag_uart_avalon_jtag_slave,
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      jtag_uart_avalon_jtag_slave_address => jtag_uart_avalon_jtag_slave_address,
      jtag_uart_avalon_jtag_slave_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      jtag_uart_avalon_jtag_slave_dataavailable_from_sa => jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      jtag_uart_avalon_jtag_slave_read_n => jtag_uart_avalon_jtag_slave_read_n,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_readyfordata_from_sa => jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
      jtag_uart_avalon_jtag_slave_reset_n => jtag_uart_avalon_jtag_slave_reset_n,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      jtag_uart_avalon_jtag_slave_write_n => jtag_uart_avalon_jtag_slave_write_n,
      jtag_uart_avalon_jtag_slave_writedata => jtag_uart_avalon_jtag_slave_writedata,
      clk => internal_pll_c2_out,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      jtag_uart_avalon_jtag_slave_dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      jtag_uart_avalon_jtag_slave_irq => jtag_uart_avalon_jtag_slave_irq,
      jtag_uart_avalon_jtag_slave_readdata => jtag_uart_avalon_jtag_slave_readdata,
      jtag_uart_avalon_jtag_slave_readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      jtag_uart_avalon_jtag_slave_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      reset_n => pll_c2_out_reset_n
    );


  --the_jtag_uart, which is an e_ptf_instance
  the_jtag_uart : jtag_uart
    port map(
      av_irq => jtag_uart_avalon_jtag_slave_irq,
      av_readdata => jtag_uart_avalon_jtag_slave_readdata,
      av_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      av_address => jtag_uart_avalon_jtag_slave_address,
      av_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      av_read_n => jtag_uart_avalon_jtag_slave_read_n,
      av_write_n => jtag_uart_avalon_jtag_slave_write_n,
      av_writedata => jtag_uart_avalon_jtag_slave_writedata,
      clk => internal_pll_c2_out,
      rst_n => jtag_uart_avalon_jtag_slave_reset_n
    );


  --the_led_pio_s1, which is an e_instance
  the_led_pio_s1 : led_pio_s1_arbitrator
    port map(
      clock_crossing_0_m1_granted_led_pio_s1 => clock_crossing_0_m1_granted_led_pio_s1,
      clock_crossing_0_m1_qualified_request_led_pio_s1 => clock_crossing_0_m1_qualified_request_led_pio_s1,
      clock_crossing_0_m1_read_data_valid_led_pio_s1 => clock_crossing_0_m1_read_data_valid_led_pio_s1,
      clock_crossing_0_m1_requests_led_pio_s1 => clock_crossing_0_m1_requests_led_pio_s1,
      d1_led_pio_s1_end_xfer => d1_led_pio_s1_end_xfer,
      led_pio_s1_address => led_pio_s1_address,
      led_pio_s1_chipselect => led_pio_s1_chipselect,
      led_pio_s1_readdata_from_sa => led_pio_s1_readdata_from_sa,
      led_pio_s1_reset_n => led_pio_s1_reset_n,
      led_pio_s1_write_n => led_pio_s1_write_n,
      led_pio_s1_writedata => led_pio_s1_writedata,
      clk => internal_pll_c2_out,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      led_pio_s1_readdata => led_pio_s1_readdata,
      reset_n => pll_c2_out_reset_n
    );


  --the_led_pio, which is an e_ptf_instance
  the_led_pio : led_pio
    port map(
      out_port => internal_out_port_from_the_led_pio,
      readdata => led_pio_s1_readdata,
      address => led_pio_s1_address,
      chipselect => led_pio_s1_chipselect,
      clk => internal_pll_c2_out,
      reset_n => led_pio_s1_reset_n,
      write_n => led_pio_s1_write_n,
      writedata => led_pio_s1_writedata
    );


  --the_onchip_memory_s1, which is an e_instance
  the_onchip_memory_s1 : onchip_memory_s1_arbitrator
    port map(
      cpu_0_data_master_granted_onchip_memory_s1 => cpu_0_data_master_granted_onchip_memory_s1,
      cpu_0_data_master_qualified_request_onchip_memory_s1 => cpu_0_data_master_qualified_request_onchip_memory_s1,
      cpu_0_data_master_read_data_valid_onchip_memory_s1 => cpu_0_data_master_read_data_valid_onchip_memory_s1,
      cpu_0_data_master_requests_onchip_memory_s1 => cpu_0_data_master_requests_onchip_memory_s1,
      cpu_0_instruction_master_granted_onchip_memory_s1 => cpu_0_instruction_master_granted_onchip_memory_s1,
      cpu_0_instruction_master_qualified_request_onchip_memory_s1 => cpu_0_instruction_master_qualified_request_onchip_memory_s1,
      cpu_0_instruction_master_read_data_valid_onchip_memory_s1 => cpu_0_instruction_master_read_data_valid_onchip_memory_s1,
      cpu_0_instruction_master_requests_onchip_memory_s1 => cpu_0_instruction_master_requests_onchip_memory_s1,
      d1_onchip_memory_s1_end_xfer => d1_onchip_memory_s1_end_xfer,
      onchip_memory_s1_address => onchip_memory_s1_address,
      onchip_memory_s1_byteenable => onchip_memory_s1_byteenable,
      onchip_memory_s1_chipselect => onchip_memory_s1_chipselect,
      onchip_memory_s1_clken => onchip_memory_s1_clken,
      onchip_memory_s1_readdata_from_sa => onchip_memory_s1_readdata_from_sa,
      onchip_memory_s1_reset => onchip_memory_s1_reset,
      onchip_memory_s1_write => onchip_memory_s1_write,
      onchip_memory_s1_writedata => onchip_memory_s1_writedata,
      registered_cpu_0_data_master_read_data_valid_onchip_memory_s1 => registered_cpu_0_data_master_read_data_valid_onchip_memory_s1,
      clk => internal_cpu_clk,
      cpu_0_data_master_address_to_slave => cpu_0_data_master_address_to_slave,
      cpu_0_data_master_byteenable => cpu_0_data_master_byteenable,
      cpu_0_data_master_read => cpu_0_data_master_read,
      cpu_0_data_master_waitrequest => cpu_0_data_master_waitrequest,
      cpu_0_data_master_write => cpu_0_data_master_write,
      cpu_0_data_master_writedata => cpu_0_data_master_writedata,
      cpu_0_instruction_master_address_to_slave => cpu_0_instruction_master_address_to_slave,
      cpu_0_instruction_master_read => cpu_0_instruction_master_read,
      onchip_memory_s1_readdata => onchip_memory_s1_readdata,
      reset_n => cpu_clk_reset_n
    );


  --the_onchip_memory, which is an e_ptf_instance
  the_onchip_memory : onchip_memory
    port map(
      readdata => onchip_memory_s1_readdata,
      address => onchip_memory_s1_address,
      byteenable => onchip_memory_s1_byteenable,
      chipselect => onchip_memory_s1_chipselect,
      clk => internal_cpu_clk,
      clken => onchip_memory_s1_clken,
      reset => onchip_memory_s1_reset,
      write => onchip_memory_s1_write,
      writedata => onchip_memory_s1_writedata
    );


  --the_pipeline_bridge_before_tristate_s1, which is an e_instance
  the_pipeline_bridge_before_tristate_s1 : pipeline_bridge_before_tristate_s1_arbitrator
    port map(
      d1_pipeline_bridge_before_tristate_s1_end_xfer => d1_pipeline_bridge_before_tristate_s1_end_xfer,
      flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1 => flash_ssram_pipeline_bridge_m1_granted_pipeline_bridge_before_tristate_s1,
      flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1 => flash_ssram_pipeline_bridge_m1_qualified_request_pipeline_bridge_before_tristate_s1,
      flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1 => flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1,
      flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1_shift_register => flash_ssram_pipeline_bridge_m1_read_data_valid_pipeline_bridge_before_tristate_s1_shift_register,
      flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1 => flash_ssram_pipeline_bridge_m1_requests_pipeline_bridge_before_tristate_s1,
      pipeline_bridge_before_tristate_s1_address => pipeline_bridge_before_tristate_s1_address,
      pipeline_bridge_before_tristate_s1_arbiterlock => pipeline_bridge_before_tristate_s1_arbiterlock,
      pipeline_bridge_before_tristate_s1_arbiterlock2 => pipeline_bridge_before_tristate_s1_arbiterlock2,
      pipeline_bridge_before_tristate_s1_burstcount => pipeline_bridge_before_tristate_s1_burstcount,
      pipeline_bridge_before_tristate_s1_byteenable => pipeline_bridge_before_tristate_s1_byteenable,
      pipeline_bridge_before_tristate_s1_chipselect => pipeline_bridge_before_tristate_s1_chipselect,
      pipeline_bridge_before_tristate_s1_debugaccess => pipeline_bridge_before_tristate_s1_debugaccess,
      pipeline_bridge_before_tristate_s1_endofpacket_from_sa => pipeline_bridge_before_tristate_s1_endofpacket_from_sa,
      pipeline_bridge_before_tristate_s1_nativeaddress => pipeline_bridge_before_tristate_s1_nativeaddress,
      pipeline_bridge_before_tristate_s1_read => pipeline_bridge_before_tristate_s1_read,
      pipeline_bridge_before_tristate_s1_readdata_from_sa => pipeline_bridge_before_tristate_s1_readdata_from_sa,
      pipeline_bridge_before_tristate_s1_reset_n => pipeline_bridge_before_tristate_s1_reset_n,
      pipeline_bridge_before_tristate_s1_waitrequest_from_sa => pipeline_bridge_before_tristate_s1_waitrequest_from_sa,
      pipeline_bridge_before_tristate_s1_write => pipeline_bridge_before_tristate_s1_write,
      pipeline_bridge_before_tristate_s1_writedata => pipeline_bridge_before_tristate_s1_writedata,
      clk => internal_cpu_clk,
      flash_ssram_pipeline_bridge_m1_address_to_slave => flash_ssram_pipeline_bridge_m1_address_to_slave,
      flash_ssram_pipeline_bridge_m1_burstcount => flash_ssram_pipeline_bridge_m1_burstcount,
      flash_ssram_pipeline_bridge_m1_byteenable => flash_ssram_pipeline_bridge_m1_byteenable,
      flash_ssram_pipeline_bridge_m1_chipselect => flash_ssram_pipeline_bridge_m1_chipselect,
      flash_ssram_pipeline_bridge_m1_debugaccess => flash_ssram_pipeline_bridge_m1_debugaccess,
      flash_ssram_pipeline_bridge_m1_latency_counter => flash_ssram_pipeline_bridge_m1_latency_counter,
      flash_ssram_pipeline_bridge_m1_read => flash_ssram_pipeline_bridge_m1_read,
      flash_ssram_pipeline_bridge_m1_write => flash_ssram_pipeline_bridge_m1_write,
      flash_ssram_pipeline_bridge_m1_writedata => flash_ssram_pipeline_bridge_m1_writedata,
      pipeline_bridge_before_tristate_s1_endofpacket => pipeline_bridge_before_tristate_s1_endofpacket,
      pipeline_bridge_before_tristate_s1_readdata => pipeline_bridge_before_tristate_s1_readdata,
      pipeline_bridge_before_tristate_s1_readdatavalid => pipeline_bridge_before_tristate_s1_readdatavalid,
      pipeline_bridge_before_tristate_s1_waitrequest => pipeline_bridge_before_tristate_s1_waitrequest,
      reset_n => cpu_clk_reset_n
    );


  --the_pipeline_bridge_before_tristate_m1, which is an e_instance
  the_pipeline_bridge_before_tristate_m1 : pipeline_bridge_before_tristate_m1_arbitrator
    port map(
      pipeline_bridge_before_tristate_m1_address_to_slave => pipeline_bridge_before_tristate_m1_address_to_slave,
      pipeline_bridge_before_tristate_m1_dbs_address => pipeline_bridge_before_tristate_m1_dbs_address,
      pipeline_bridge_before_tristate_m1_dbs_write_16 => pipeline_bridge_before_tristate_m1_dbs_write_16,
      pipeline_bridge_before_tristate_m1_latency_counter => pipeline_bridge_before_tristate_m1_latency_counter,
      pipeline_bridge_before_tristate_m1_readdata => pipeline_bridge_before_tristate_m1_readdata,
      pipeline_bridge_before_tristate_m1_readdatavalid => pipeline_bridge_before_tristate_m1_readdatavalid,
      pipeline_bridge_before_tristate_m1_waitrequest => pipeline_bridge_before_tristate_m1_waitrequest,
      cfi_flash_s1_wait_counter_eq_0 => cfi_flash_s1_wait_counter_eq_0,
      clk => internal_cpu_clk,
      d1_flash_ssram_tristate_avalon_slave_end_xfer => d1_flash_ssram_tristate_avalon_slave_end_xfer,
      incoming_flash_ssram_tristate_data => incoming_flash_ssram_tristate_data,
      incoming_flash_ssram_tristate_data_with_Xs_converted_to_0 => incoming_flash_ssram_tristate_data_with_Xs_converted_to_0,
      pipeline_bridge_before_tristate_m1_address => pipeline_bridge_before_tristate_m1_address,
      pipeline_bridge_before_tristate_m1_burstcount => pipeline_bridge_before_tristate_m1_burstcount,
      pipeline_bridge_before_tristate_m1_byteenable => pipeline_bridge_before_tristate_m1_byteenable,
      pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1 => pipeline_bridge_before_tristate_m1_byteenable_cfi_flash_s1,
      pipeline_bridge_before_tristate_m1_chipselect => pipeline_bridge_before_tristate_m1_chipselect,
      pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1 => pipeline_bridge_before_tristate_m1_granted_cfi_flash_s1,
      pipeline_bridge_before_tristate_m1_granted_ssram_s1 => pipeline_bridge_before_tristate_m1_granted_ssram_s1,
      pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1 => pipeline_bridge_before_tristate_m1_qualified_request_cfi_flash_s1,
      pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1 => pipeline_bridge_before_tristate_m1_qualified_request_ssram_s1,
      pipeline_bridge_before_tristate_m1_read => pipeline_bridge_before_tristate_m1_read,
      pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1 => pipeline_bridge_before_tristate_m1_read_data_valid_cfi_flash_s1,
      pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1 => pipeline_bridge_before_tristate_m1_read_data_valid_ssram_s1,
      pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1 => pipeline_bridge_before_tristate_m1_requests_cfi_flash_s1,
      pipeline_bridge_before_tristate_m1_requests_ssram_s1 => pipeline_bridge_before_tristate_m1_requests_ssram_s1,
      pipeline_bridge_before_tristate_m1_write => pipeline_bridge_before_tristate_m1_write,
      pipeline_bridge_before_tristate_m1_writedata => pipeline_bridge_before_tristate_m1_writedata,
      reset_n => cpu_clk_reset_n
    );


  --the_pipeline_bridge_before_tristate, which is an e_ptf_instance
  the_pipeline_bridge_before_tristate : pipeline_bridge_before_tristate
    port map(
      m1_address => pipeline_bridge_before_tristate_m1_address,
      m1_burstcount => pipeline_bridge_before_tristate_m1_burstcount,
      m1_byteenable => pipeline_bridge_before_tristate_m1_byteenable,
      m1_chipselect => pipeline_bridge_before_tristate_m1_chipselect,
      m1_debugaccess => pipeline_bridge_before_tristate_m1_debugaccess,
      m1_read => pipeline_bridge_before_tristate_m1_read,
      m1_write => pipeline_bridge_before_tristate_m1_write,
      m1_writedata => pipeline_bridge_before_tristate_m1_writedata,
      s1_endofpacket => pipeline_bridge_before_tristate_s1_endofpacket,
      s1_readdata => pipeline_bridge_before_tristate_s1_readdata,
      s1_readdatavalid => pipeline_bridge_before_tristate_s1_readdatavalid,
      s1_waitrequest => pipeline_bridge_before_tristate_s1_waitrequest,
      clk => internal_cpu_clk,
      m1_endofpacket => pipeline_bridge_before_tristate_m1_endofpacket,
      m1_readdata => pipeline_bridge_before_tristate_m1_readdata,
      m1_readdatavalid => pipeline_bridge_before_tristate_m1_readdatavalid,
      m1_waitrequest => pipeline_bridge_before_tristate_m1_waitrequest,
      reset_n => pipeline_bridge_before_tristate_s1_reset_n,
      s1_address => pipeline_bridge_before_tristate_s1_address,
      s1_arbiterlock => pipeline_bridge_before_tristate_s1_arbiterlock,
      s1_arbiterlock2 => pipeline_bridge_before_tristate_s1_arbiterlock2,
      s1_burstcount => pipeline_bridge_before_tristate_s1_burstcount,
      s1_byteenable => pipeline_bridge_before_tristate_s1_byteenable,
      s1_chipselect => pipeline_bridge_before_tristate_s1_chipselect,
      s1_debugaccess => pipeline_bridge_before_tristate_s1_debugaccess,
      s1_nativeaddress => pipeline_bridge_before_tristate_s1_nativeaddress,
      s1_read => pipeline_bridge_before_tristate_s1_read,
      s1_write => pipeline_bridge_before_tristate_s1_write,
      s1_writedata => pipeline_bridge_before_tristate_s1_writedata
    );


  --the_pll_s1, which is an e_instance
  the_pll_s1 : pll_s1_arbitrator
    port map(
      d1_pll_s1_end_xfer => d1_pll_s1_end_xfer,
      gpib_edm1_clock_0_out_granted_pll_s1 => gpib_edm1_clock_0_out_granted_pll_s1,
      gpib_edm1_clock_0_out_qualified_request_pll_s1 => gpib_edm1_clock_0_out_qualified_request_pll_s1,
      gpib_edm1_clock_0_out_read_data_valid_pll_s1 => gpib_edm1_clock_0_out_read_data_valid_pll_s1,
      gpib_edm1_clock_0_out_requests_pll_s1 => gpib_edm1_clock_0_out_requests_pll_s1,
      pll_s1_address => pll_s1_address,
      pll_s1_chipselect => pll_s1_chipselect,
      pll_s1_read => pll_s1_read,
      pll_s1_readdata_from_sa => pll_s1_readdata_from_sa,
      pll_s1_reset_n => pll_s1_reset_n,
      pll_s1_resetrequest_from_sa => pll_s1_resetrequest_from_sa,
      pll_s1_write => pll_s1_write,
      pll_s1_writedata => pll_s1_writedata,
      clk => clk_0,
      gpib_edm1_clock_0_out_address_to_slave => gpib_edm1_clock_0_out_address_to_slave,
      gpib_edm1_clock_0_out_nativeaddress => gpib_edm1_clock_0_out_nativeaddress,
      gpib_edm1_clock_0_out_read => gpib_edm1_clock_0_out_read,
      gpib_edm1_clock_0_out_write => gpib_edm1_clock_0_out_write,
      gpib_edm1_clock_0_out_writedata => gpib_edm1_clock_0_out_writedata,
      pll_s1_readdata => pll_s1_readdata,
      pll_s1_resetrequest => pll_s1_resetrequest,
      reset_n => clk_0_reset_n
    );


  --cpu_clk out_clk assignment, which is an e_assign
  internal_cpu_clk <= out_clk_pll_c0;
  --ssram_clk out_clk assignment, which is an e_assign
  ssram_clk <= out_clk_pll_c1;
  --pll_c2_out out_clk assignment, which is an e_assign
  internal_pll_c2_out <= out_clk_pll_c2;
  --pll_c3_out out_clk assignment, which is an e_assign
  internal_pll_c3_out <= out_clk_pll_c3;
  --the_pll, which is an e_ptf_instance
  the_pll : pll
    port map(
      c0 => out_clk_pll_c0,
      c1 => out_clk_pll_c1,
      c2 => out_clk_pll_c2,
      c3 => out_clk_pll_c3,
      readdata => pll_s1_readdata,
      resetrequest => pll_s1_resetrequest,
      address => pll_s1_address,
      chipselect => pll_s1_chipselect,
      clk => clk_0,
      read => pll_s1_read,
      reset_n => pll_s1_reset_n,
      write => pll_s1_write,
      writedata => pll_s1_writedata
    );


  --the_remote_update_cycloneiii_1_s1, which is an e_instance
  the_remote_update_cycloneiii_1_s1 : remote_update_cycloneiii_1_s1_arbitrator
    port map(
      d1_remote_update_cycloneiii_1_s1_end_xfer => d1_remote_update_cycloneiii_1_s1_end_xfer,
      gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1 => gpib_edm1_clock_1_out_granted_remote_update_cycloneiii_1_s1,
      gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1 => gpib_edm1_clock_1_out_qualified_request_remote_update_cycloneiii_1_s1,
      gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1 => gpib_edm1_clock_1_out_read_data_valid_remote_update_cycloneiii_1_s1,
      gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1 => gpib_edm1_clock_1_out_requests_remote_update_cycloneiii_1_s1,
      remote_update_cycloneiii_1_s1_address => remote_update_cycloneiii_1_s1_address,
      remote_update_cycloneiii_1_s1_chipselect => remote_update_cycloneiii_1_s1_chipselect,
      remote_update_cycloneiii_1_s1_read => remote_update_cycloneiii_1_s1_read,
      remote_update_cycloneiii_1_s1_readdata_from_sa => remote_update_cycloneiii_1_s1_readdata_from_sa,
      remote_update_cycloneiii_1_s1_reset => remote_update_cycloneiii_1_s1_reset,
      remote_update_cycloneiii_1_s1_waitrequest_from_sa => remote_update_cycloneiii_1_s1_waitrequest_from_sa,
      remote_update_cycloneiii_1_s1_write => remote_update_cycloneiii_1_s1_write,
      remote_update_cycloneiii_1_s1_writedata => remote_update_cycloneiii_1_s1_writedata,
      clk => internal_pll_c3_out,
      gpib_edm1_clock_1_out_address_to_slave => gpib_edm1_clock_1_out_address_to_slave,
      gpib_edm1_clock_1_out_nativeaddress => gpib_edm1_clock_1_out_nativeaddress,
      gpib_edm1_clock_1_out_read => gpib_edm1_clock_1_out_read,
      gpib_edm1_clock_1_out_write => gpib_edm1_clock_1_out_write,
      gpib_edm1_clock_1_out_writedata => gpib_edm1_clock_1_out_writedata,
      remote_update_cycloneiii_1_s1_readdata => remote_update_cycloneiii_1_s1_readdata,
      remote_update_cycloneiii_1_s1_waitrequest => remote_update_cycloneiii_1_s1_waitrequest,
      reset_n => pll_c3_out_reset_n
    );


  --the_remote_update_cycloneiii_1, which is an e_ptf_instance
  the_remote_update_cycloneiii_1 : remote_update_cycloneiii_1
    port map(
      readdata => remote_update_cycloneiii_1_s1_readdata,
      waitrequest => remote_update_cycloneiii_1_s1_waitrequest,
      address => remote_update_cycloneiii_1_s1_address,
      chipselect => remote_update_cycloneiii_1_s1_chipselect,
      clk => internal_pll_c3_out,
      read => remote_update_cycloneiii_1_s1_read,
      reset => remote_update_cycloneiii_1_s1_reset,
      write => remote_update_cycloneiii_1_s1_write,
      writedata => remote_update_cycloneiii_1_s1_writedata
    );


  --the_sys_clk_s1, which is an e_instance
  the_sys_clk_s1 : sys_clk_s1_arbitrator
    port map(
      clock_crossing_0_m1_granted_sys_clk_s1 => clock_crossing_0_m1_granted_sys_clk_s1,
      clock_crossing_0_m1_qualified_request_sys_clk_s1 => clock_crossing_0_m1_qualified_request_sys_clk_s1,
      clock_crossing_0_m1_read_data_valid_sys_clk_s1 => clock_crossing_0_m1_read_data_valid_sys_clk_s1,
      clock_crossing_0_m1_requests_sys_clk_s1 => clock_crossing_0_m1_requests_sys_clk_s1,
      d1_sys_clk_s1_end_xfer => d1_sys_clk_s1_end_xfer,
      sys_clk_s1_address => sys_clk_s1_address,
      sys_clk_s1_chipselect => sys_clk_s1_chipselect,
      sys_clk_s1_irq_from_sa => sys_clk_s1_irq_from_sa,
      sys_clk_s1_readdata_from_sa => sys_clk_s1_readdata_from_sa,
      sys_clk_s1_reset_n => sys_clk_s1_reset_n,
      sys_clk_s1_write_n => sys_clk_s1_write_n,
      sys_clk_s1_writedata => sys_clk_s1_writedata,
      clk => internal_pll_c2_out,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      reset_n => pll_c2_out_reset_n,
      sys_clk_s1_irq => sys_clk_s1_irq,
      sys_clk_s1_readdata => sys_clk_s1_readdata
    );


  --the_sys_clk, which is an e_ptf_instance
  the_sys_clk : sys_clk
    port map(
      irq => sys_clk_s1_irq,
      readdata => sys_clk_s1_readdata,
      address => sys_clk_s1_address,
      chipselect => sys_clk_s1_chipselect,
      clk => internal_pll_c2_out,
      reset_n => sys_clk_s1_reset_n,
      write_n => sys_clk_s1_write_n,
      writedata => sys_clk_s1_writedata
    );


  --reset is asserted asynchronously and deasserted synchronously
  gpib_edm1_reset_cpu_clk_domain_synch : gpib_edm1_reset_cpu_clk_domain_synch_module
    port map(
      data_out => cpu_clk_reset_n,
      clk => internal_cpu_clk,
      data_in => module_input25,
      reset_n => reset_n_sources
    );

  module_input25 <= std_logic'('1');

  --reset is asserted asynchronously and deasserted synchronously
  gpib_edm1_reset_ddr_sdram_phy_clk_out_domain_synch : gpib_edm1_reset_ddr_sdram_phy_clk_out_domain_synch_module
    port map(
      data_out => ddr_sdram_phy_clk_out_reset_n,
      clk => internal_ddr_sdram_phy_clk_out,
      data_in => module_input26,
      reset_n => reset_n_sources
    );

  module_input26 <= std_logic'('1');

  --reset is asserted asynchronously and deasserted synchronously
  gpib_edm1_reset_pll_c2_out_domain_synch : gpib_edm1_reset_pll_c2_out_domain_synch_module
    port map(
      data_out => pll_c2_out_reset_n,
      clk => internal_pll_c2_out,
      data_in => module_input27,
      reset_n => reset_n_sources
    );

  module_input27 <= std_logic'('1');

  --reset is asserted asynchronously and deasserted synchronously
  gpib_edm1_reset_pll_c3_out_domain_synch : gpib_edm1_reset_pll_c3_out_domain_synch_module
    port map(
      data_out => pll_c3_out_reset_n,
      clk => internal_pll_c3_out,
      data_in => module_input28,
      reset_n => reset_n_sources
    );

  module_input28 <= std_logic'('1');

  --cpu_ddr_clock_bridge_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  cpu_ddr_clock_bridge_m1_endofpacket <= std_logic'('0');
  --gpib_edm1_clock_0_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  gpib_edm1_clock_0_out_endofpacket <= std_logic'('0');
  --gpib_edm1_clock_1_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  gpib_edm1_clock_1_out_endofpacket <= std_logic'('0');
  --pipeline_bridge_before_tristate_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  pipeline_bridge_before_tristate_m1_endofpacket <= std_logic'('0');
  --vhdl renameroo for output signals
  MOSI_from_the_ad7928 <= internal_MOSI_from_the_ad7928;
  --vhdl renameroo for output signals
  MOSI_from_the_dac_ad5308 <= internal_MOSI_from_the_dac_ad5308;
  --vhdl renameroo for output signals
  SCLK_from_the_ad7928 <= internal_SCLK_from_the_ad7928;
  --vhdl renameroo for output signals
  SCLK_from_the_dac_ad5308 <= internal_SCLK_from_the_dac_ad5308;
  --vhdl renameroo for output signals
  SS_n_from_the_ad7928 <= internal_SS_n_from_the_ad7928;
  --vhdl renameroo for output signals
  SS_n_from_the_dac_ad5308 <= internal_SS_n_from_the_dac_ad5308;
  --vhdl renameroo for output signals
  adsc_n_to_the_ssram <= internal_adsc_n_to_the_ssram;
  --vhdl renameroo for output signals
  bw_n_to_the_ssram <= internal_bw_n_to_the_ssram;
  --vhdl renameroo for output signals
  bwe_n_to_the_ssram <= internal_bwe_n_to_the_ssram;
  --vhdl renameroo for output signals
  chipenable1_n_to_the_ssram <= internal_chipenable1_n_to_the_ssram;
  --vhdl renameroo for output signals
  cpu_clk <= internal_cpu_clk;
  --vhdl renameroo for output signals
  ddr_sdram_phy_clk_out <= internal_ddr_sdram_phy_clk_out;
  --vhdl renameroo for output signals
  flash_ssram_tristate_address <= internal_flash_ssram_tristate_address;
  --vhdl renameroo for output signals
  local_init_done_from_the_ddr_sdram <= internal_local_init_done_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  local_refresh_ack_from_the_ddr_sdram <= internal_local_refresh_ack_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  local_wdata_req_from_the_ddr_sdram <= internal_local_wdata_req_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  mem_addr_from_the_ddr_sdram <= internal_mem_addr_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  mem_ba_from_the_ddr_sdram <= internal_mem_ba_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  mem_cas_n_from_the_ddr_sdram <= internal_mem_cas_n_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  mem_cke_from_the_ddr_sdram <= internal_mem_cke_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  mem_cs_n_from_the_ddr_sdram <= internal_mem_cs_n_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  mem_dm_from_the_ddr_sdram <= internal_mem_dm_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  mem_ras_n_from_the_ddr_sdram <= internal_mem_ras_n_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  mem_we_n_from_the_ddr_sdram <= internal_mem_we_n_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  out_port_from_the_gpib_leds <= internal_out_port_from_the_gpib_leds;
  --vhdl renameroo for output signals
  out_port_from_the_gpio2 <= internal_out_port_from_the_gpio2;
  --vhdl renameroo for output signals
  out_port_from_the_led_pio <= internal_out_port_from_the_led_pio;
  --vhdl renameroo for output signals
  outputenable_n_to_the_ssram <= internal_outputenable_n_to_the_ssram;
  --vhdl renameroo for output signals
  pll_c2_out <= internal_pll_c2_out;
  --vhdl renameroo for output signals
  pll_c3_out <= internal_pll_c3_out;
  --vhdl renameroo for output signals
  read_n_to_the_cfi_flash <= internal_read_n_to_the_cfi_flash;
  --vhdl renameroo for output signals
  reset_n_to_the_ssram <= internal_reset_n_to_the_ssram;
  --vhdl renameroo for output signals
  reset_phy_clk_n_from_the_ddr_sdram <= internal_reset_phy_clk_n_from_the_ddr_sdram;
  --vhdl renameroo for output signals
  select_n_to_the_cfi_flash <= internal_select_n_to_the_cfi_flash;
  --vhdl renameroo for output signals
  write_n_to_the_cfi_flash <= internal_write_n_to_the_cfi_flash;

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cfi_flash_lane0_module is 
        port (
              -- inputs:
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity cfi_flash_lane0_module;


architecture europa of cfi_flash_lane0_module is
              signal internal_q :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 8388607 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, rdaddress) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (22 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "cfi_flash_lane0.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 8388608) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rdaddress)));
      


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity cfi_flash_lane0_module is 
--        port (
--              
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity cfi_flash_lane0_module;
--
--
--architecture europa of cfi_flash_lane0_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal internal_q :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 8388607 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
--
--begin
--
--  process (rdaddress)
--  begin
--      read_address <= rdaddress;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "cfi_flash_lane0.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "UNREGISTERED",
--      lpm_rdaddress_control => "UNREGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 23,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cfi_flash_lane1_module is 
        port (
              -- inputs:
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity cfi_flash_lane1_module;


architecture europa of cfi_flash_lane1_module is
              signal internal_q1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 8388607 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, rdaddress) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (22 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "cfi_flash_lane1.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 8388608) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rdaddress)));
      


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity cfi_flash_lane1_module is 
--        port (
--              
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity cfi_flash_lane1_module;
--
--
--architecture europa of cfi_flash_lane1_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal internal_q1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 8388607 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
--
--begin
--
--  process (rdaddress)
--  begin
--      read_address <= rdaddress;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "cfi_flash_lane1.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "UNREGISTERED",
--      lpm_rdaddress_control => "UNREGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 23,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q1,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q1;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cfi_flash is 
        port (
              -- inputs:
                 signal address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal read_n : IN STD_LOGIC;
                 signal select_n : IN STD_LOGIC;
                 signal write_n : IN STD_LOGIC;

              -- outputs:
                 signal data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity cfi_flash;


architecture europa of cfi_flash is
--synthesis translate_off
component cfi_flash_lane0_module is 
           port (
                 -- inputs:
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component cfi_flash_lane0_module;

component cfi_flash_lane1_module is 
           port (
                 -- inputs:
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component cfi_flash_lane1_module;

--synthesis translate_on
                signal data_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal data_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal logic_vector_gasket :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal module_input29 :  STD_LOGIC;
                signal module_input30 :  STD_LOGIC;
                signal module_input31 :  STD_LOGIC;
                signal module_input32 :  STD_LOGIC;
                signal q_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal q_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);

begin

  --s1, which is an e_ptf_slave
--synthesis translate_off
    logic_vector_gasket <= data;
    data_0 <= logic_vector_gasket(7 DOWNTO 0);
    --cfi_flash_lane0, which is an e_ram
    cfi_flash_lane0 : cfi_flash_lane0_module
      port map(
        q => q_0,
        data => data_0,
        rdaddress => address,
        rdclken => module_input29,
        wraddress => address,
        wrclock => write_n,
        wren => module_input30
      );

    module_input29 <= std_logic'('1');
    module_input30 <= NOT select_n;

    data_1 <= logic_vector_gasket(15 DOWNTO 8);
    --cfi_flash_lane1, which is an e_ram
    cfi_flash_lane1 : cfi_flash_lane1_module
      port map(
        q => q_1,
        data => data_1,
        rdaddress => address,
        rdclken => module_input31,
        wraddress => address,
        wrclock => write_n,
        wren => module_input32
      );

    module_input31 <= std_logic'('1');
    module_input32 <= NOT select_n;

    data <= A_WE_StdLogicVector((std_logic'(((NOT select_n AND NOT read_n))) = '1'), (q_1 & q_0), A_REP(std_logic'('Z'), 16));
--synthesis translate_on

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ssram_lane0_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ssram_lane0_module;


architecture europa of ssram_lane0_module is
              signal d1_rdaddress :  STD_LOGIC_VECTOR (17 DOWNTO 0);
              signal internal_q2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 262143 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, clk) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;
    VARIABLE rd_address_internal : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');
    VARIABLE d1_rdaddress : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "ssram_lane0.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 262144) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rd_address_internal)));
      
			 IF clk'event AND clk = '1' AND rdclken = '1' THEN
                            rd_address_internal := d1_rdaddress;
                            d1_rdaddress := rdaddress;

                         END IF;
                        


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity ssram_lane0_module is 
--        port (
--              
--                 signal clk : IN STD_LOGIC;
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal reset_n : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity ssram_lane0_module;
--
--
--architecture europa of ssram_lane0_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal rdclock : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal d1_rdaddress :  STD_LOGIC_VECTOR (17 DOWNTO 0);
--                signal internal_q2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 262143 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);
--
--begin
--
--  process (rdaddress)
--  begin
--      read_address <= rdaddress;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "ssram_lane0.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "REGISTERED",
--      lpm_rdaddress_control => "REGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 18,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q2,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            rdclock => clk,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q2;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ssram_lane1_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ssram_lane1_module;


architecture europa of ssram_lane1_module is
              signal d1_rdaddress :  STD_LOGIC_VECTOR (17 DOWNTO 0);
              signal internal_q3 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 262143 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, clk) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;
    VARIABLE rd_address_internal : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');
    VARIABLE d1_rdaddress : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "ssram_lane1.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 262144) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rd_address_internal)));
      
			 IF clk'event AND clk = '1' AND rdclken = '1' THEN
                            rd_address_internal := d1_rdaddress;
                            d1_rdaddress := rdaddress;

                         END IF;
                        


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity ssram_lane1_module is 
--        port (
--              
--                 signal clk : IN STD_LOGIC;
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal reset_n : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity ssram_lane1_module;
--
--
--architecture europa of ssram_lane1_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal rdclock : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal d1_rdaddress :  STD_LOGIC_VECTOR (17 DOWNTO 0);
--                signal internal_q3 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 262143 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);
--
--begin
--
--  process (rdaddress)
--  begin
--      read_address <= rdaddress;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "ssram_lane1.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "REGISTERED",
--      lpm_rdaddress_control => "REGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 18,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q3,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            rdclock => clk,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q3;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ssram_lane2_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ssram_lane2_module;


architecture europa of ssram_lane2_module is
              signal d1_rdaddress :  STD_LOGIC_VECTOR (17 DOWNTO 0);
              signal internal_q4 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 262143 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, clk) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;
    VARIABLE rd_address_internal : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');
    VARIABLE d1_rdaddress : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "ssram_lane2.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 262144) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rd_address_internal)));
      
			 IF clk'event AND clk = '1' AND rdclken = '1' THEN
                            rd_address_internal := d1_rdaddress;
                            d1_rdaddress := rdaddress;

                         END IF;
                        


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity ssram_lane2_module is 
--        port (
--              
--                 signal clk : IN STD_LOGIC;
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal reset_n : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity ssram_lane2_module;
--
--
--architecture europa of ssram_lane2_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal rdclock : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal d1_rdaddress :  STD_LOGIC_VECTOR (17 DOWNTO 0);
--                signal internal_q4 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 262143 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);
--
--begin
--
--  process (rdaddress)
--  begin
--      read_address <= rdaddress;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "ssram_lane2.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "REGISTERED",
--      lpm_rdaddress_control => "REGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 18,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q4,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            rdclock => clk,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q4;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ssram_lane3_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ssram_lane3_module;


architecture europa of ssram_lane3_module is
              signal d1_rdaddress :  STD_LOGIC_VECTOR (17 DOWNTO 0);
              signal internal_q5 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 262143 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, clk) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;
    VARIABLE rd_address_internal : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');
    VARIABLE d1_rdaddress : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (17 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "ssram_lane3.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 262144) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rd_address_internal)));
      
			 IF clk'event AND clk = '1' AND rdclken = '1' THEN
                            rd_address_internal := d1_rdaddress;
                            d1_rdaddress := rdaddress;

                         END IF;
                        


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity ssram_lane3_module is 
--        port (
--              
--                 signal clk : IN STD_LOGIC;
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal reset_n : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity ssram_lane3_module;
--
--
--architecture europa of ssram_lane3_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal rdclock : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal d1_rdaddress :  STD_LOGIC_VECTOR (17 DOWNTO 0);
--                signal internal_q5 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 262143 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (17 DOWNTO 0);
--
--begin
--
--  process (rdaddress)
--  begin
--      read_address <= rdaddress;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "ssram_lane3.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "REGISTERED",
--      lpm_rdaddress_control => "REGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 18,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q5,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            rdclock => clk,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q5;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ssram is 
        port (
              -- inputs:
                 signal address : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal adsc_n : IN STD_LOGIC;
                 signal bw_n : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal bwe_n : IN STD_LOGIC;
                 signal chipenable1_n : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal outputenable_n : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity ssram;


architecture europa of ssram is
--synthesis translate_off
component ssram_lane0_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ssram_lane0_module;

component ssram_lane1_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ssram_lane1_module;

component ssram_lane2_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ssram_lane2_module;

component ssram_lane3_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ssram_lane3_module;

--synthesis translate_on
                signal data_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal data_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal data_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal data_3 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal logic_vector_gasket :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal module_input34 :  STD_LOGIC;
                signal module_input35 :  STD_LOGIC;
                signal module_input36 :  STD_LOGIC;
                signal module_input37 :  STD_LOGIC;
                signal module_input38 :  STD_LOGIC;
                signal module_input39 :  STD_LOGIC;
                signal module_input40 :  STD_LOGIC;
                signal module_input41 :  STD_LOGIC;
                signal q_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal q_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal q_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal q_3 :  STD_LOGIC_VECTOR (7 DOWNTO 0);

begin

  --s1, which is an e_ptf_slave
--synthesis translate_off
    logic_vector_gasket <= data;
    data_0 <= logic_vector_gasket(7 DOWNTO 0);
    --ssram_lane0, which is an e_ram
    ssram_lane0 : ssram_lane0_module
      port map(
        q => q_0,
        clk => clk,
        data => data_0,
        rdaddress => address,
        rdclken => module_input34,
        reset_n => reset_n,
        wraddress => address,
        wrclock => clk,
        wren => module_input35
      );

    module_input34 <= std_logic'('1');
    module_input35 <= (NOT chipenable1_n AND NOT bwe_n) AND NOT bw_n(0);

    data_1 <= logic_vector_gasket(15 DOWNTO 8);
    --ssram_lane1, which is an e_ram
    ssram_lane1 : ssram_lane1_module
      port map(
        q => q_1,
        clk => clk,
        data => data_1,
        rdaddress => address,
        rdclken => module_input36,
        reset_n => reset_n,
        wraddress => address,
        wrclock => clk,
        wren => module_input37
      );

    module_input36 <= std_logic'('1');
    module_input37 <= (NOT chipenable1_n AND NOT bwe_n) AND NOT bw_n(1);

    data_2 <= logic_vector_gasket(23 DOWNTO 16);
    --ssram_lane2, which is an e_ram
    ssram_lane2 : ssram_lane2_module
      port map(
        q => q_2,
        clk => clk,
        data => data_2,
        rdaddress => address,
        rdclken => module_input38,
        reset_n => reset_n,
        wraddress => address,
        wrclock => clk,
        wren => module_input39
      );

    module_input38 <= std_logic'('1');
    module_input39 <= (NOT chipenable1_n AND NOT bwe_n) AND NOT bw_n(2);

    data_3 <= logic_vector_gasket(31 DOWNTO 24);
    --ssram_lane3, which is an e_ram
    ssram_lane3 : ssram_lane3_module
      port map(
        q => q_3,
        clk => clk,
        data => data_3,
        rdaddress => address,
        rdclken => module_input40,
        reset_n => reset_n,
        wraddress => address,
        wrclock => clk,
        wren => module_input41
      );

    module_input40 <= std_logic'('1');
    module_input41 <= (NOT chipenable1_n AND NOT bwe_n) AND NOT bw_n(3);

    data <= A_WE_StdLogicVector((std_logic'(((NOT chipenable1_n AND NOT outputenable_n))) = '1'), (q_3 & q_2 & q_1 & q_0), A_REP(std_logic'('Z'), 32));
--synthesis translate_on

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your libraries here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>

entity test_bench is 
end entity test_bench;


architecture europa of test_bench is
component gpib_edm1 is 
           port (
                 -- 1) global signals:
                    signal clk_0 : IN STD_LOGIC;
                    signal cpu_clk : OUT STD_LOGIC;
                    signal ddr_sdram_aux_full_rate_clk_out : OUT STD_LOGIC;
                    signal ddr_sdram_aux_half_rate_clk_out : OUT STD_LOGIC;
                    signal ddr_sdram_phy_clk_out : OUT STD_LOGIC;
                    signal pll_c2_out : OUT STD_LOGIC;
                    signal pll_c3_out : OUT STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal ssram_clk : OUT STD_LOGIC;

                 -- the_ad7928
                    signal MISO_to_the_ad7928 : IN STD_LOGIC;
                    signal MOSI_from_the_ad7928 : OUT STD_LOGIC;
                    signal SCLK_from_the_ad7928 : OUT STD_LOGIC;
                    signal SS_n_from_the_ad7928 : OUT STD_LOGIC;

                 -- the_dac_ad5308
                    signal MISO_to_the_dac_ad5308 : IN STD_LOGIC;
                    signal MOSI_from_the_dac_ad5308 : OUT STD_LOGIC;
                    signal SCLK_from_the_dac_ad5308 : OUT STD_LOGIC;
                    signal SS_n_from_the_dac_ad5308 : OUT STD_LOGIC;

                 -- the_ddr_sdram
                    signal global_reset_n_to_the_ddr_sdram : IN STD_LOGIC;
                    signal local_init_done_from_the_ddr_sdram : OUT STD_LOGIC;
                    signal local_refresh_ack_from_the_ddr_sdram : OUT STD_LOGIC;
                    signal local_wdata_req_from_the_ddr_sdram : OUT STD_LOGIC;
                    signal mem_addr_from_the_ddr_sdram : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal mem_ba_from_the_ddr_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_cas_n_from_the_ddr_sdram : OUT STD_LOGIC;
                    signal mem_cke_from_the_ddr_sdram : OUT STD_LOGIC;
                    signal mem_clk_n_to_and_from_the_ddr_sdram : INOUT STD_LOGIC;
                    signal mem_clk_to_and_from_the_ddr_sdram : INOUT STD_LOGIC;
                    signal mem_cs_n_from_the_ddr_sdram : OUT STD_LOGIC;
                    signal mem_dm_from_the_ddr_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_dq_to_and_from_the_ddr_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal mem_dqs_to_and_from_the_ddr_sdram : INOUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_ras_n_from_the_ddr_sdram : OUT STD_LOGIC;
                    signal mem_we_n_from_the_ddr_sdram : OUT STD_LOGIC;
                    signal reset_phy_clk_n_from_the_ddr_sdram : OUT STD_LOGIC;

                 -- the_flash_ssram_tristate_avalon_slave
                    signal adsc_n_to_the_ssram : OUT STD_LOGIC;
                    signal bw_n_to_the_ssram : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal bwe_n_to_the_ssram : OUT STD_LOGIC;
                    signal chipenable1_n_to_the_ssram : OUT STD_LOGIC;
                    signal flash_ssram_tristate_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal flash_ssram_tristate_data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal outputenable_n_to_the_ssram : OUT STD_LOGIC;
                    signal read_n_to_the_cfi_flash : OUT STD_LOGIC;
                    signal reset_n_to_the_ssram : OUT STD_LOGIC;
                    signal select_n_to_the_cfi_flash : OUT STD_LOGIC;
                    signal write_n_to_the_cfi_flash : OUT STD_LOGIC;

                 -- the_gpib_leds
                    signal out_port_from_the_gpib_leds : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_gpio1
                    signal bidir_port_to_and_from_the_gpio1 : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_gpio2
                    signal out_port_from_the_gpio2 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_led_pio
                    signal out_port_from_the_led_pio : OUT STD_LOGIC
                 );
end component gpib_edm1;

component cfi_flash is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal read_n : IN STD_LOGIC;
                    signal select_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;

                 -- outputs:
                    signal data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component cfi_flash;

component ssram is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal adsc_n : IN STD_LOGIC;
                    signal bw_n : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal bwe_n : IN STD_LOGIC;
                    signal chipenable1_n : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal outputenable_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component ssram;

                signal MISO_to_the_ad7928 :  STD_LOGIC;
                signal MISO_to_the_dac_ad5308 :  STD_LOGIC;
                signal MOSI_from_the_ad7928 :  STD_LOGIC;
                signal MOSI_from_the_dac_ad5308 :  STD_LOGIC;
                signal SCLK_from_the_ad7928 :  STD_LOGIC;
                signal SCLK_from_the_dac_ad5308 :  STD_LOGIC;
                signal SS_n_from_the_ad7928 :  STD_LOGIC;
                signal SS_n_from_the_dac_ad5308 :  STD_LOGIC;
                signal ad7928_spi_control_port_dataavailable_from_sa :  STD_LOGIC;
                signal ad7928_spi_control_port_readyfordata_from_sa :  STD_LOGIC;
                signal adsc_n_to_the_ssram :  STD_LOGIC;
                signal bidir_port_to_and_from_the_gpio1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal bw_n_to_the_ssram :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal bwe_n_to_the_ssram :  STD_LOGIC;
                signal chipenable1_n_to_the_ssram :  STD_LOGIC;
                signal clk :  STD_LOGIC;
                signal clk_0 :  STD_LOGIC;
                signal clock_crossing_0_s1_endofpacket_from_sa :  STD_LOGIC;
                signal cpu_clk :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_endofpacket :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_dataavailable_from_sa :  STD_LOGIC;
                signal dac_ad5308_spi_control_port_readyfordata_from_sa :  STD_LOGIC;
                signal ddr_sdram_aux_full_rate_clk_out :  STD_LOGIC;
                signal ddr_sdram_aux_half_rate_clk_out :  STD_LOGIC;
                signal ddr_sdram_phy_clk_out :  STD_LOGIC;
                signal flash_ssram_pipeline_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal flash_ssram_tristate_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal flash_ssram_tristate_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal global_reset_n_to_the_ddr_sdram :  STD_LOGIC;
                signal gpib_edm1_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal gpib_edm1_clock_0_out_endofpacket :  STD_LOGIC;
                signal gpib_edm1_clock_1_in_endofpacket_from_sa :  STD_LOGIC;
                signal gpib_edm1_clock_1_out_endofpacket :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal local_init_done_from_the_ddr_sdram :  STD_LOGIC;
                signal local_refresh_ack_from_the_ddr_sdram :  STD_LOGIC;
                signal local_wdata_req_from_the_ddr_sdram :  STD_LOGIC;
                signal mem_addr_from_the_ddr_sdram :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal mem_ba_from_the_ddr_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal mem_cas_n_from_the_ddr_sdram :  STD_LOGIC;
                signal mem_cke_from_the_ddr_sdram :  STD_LOGIC;
                signal mem_clk_n_to_and_from_the_ddr_sdram :  STD_LOGIC;
                signal mem_clk_to_and_from_the_ddr_sdram :  STD_LOGIC;
                signal mem_cs_n_from_the_ddr_sdram :  STD_LOGIC;
                signal mem_dm_from_the_ddr_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal mem_dq_to_and_from_the_ddr_sdram :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal mem_dqs_to_and_from_the_ddr_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal mem_ras_n_from_the_ddr_sdram :  STD_LOGIC;
                signal mem_we_n_from_the_ddr_sdram :  STD_LOGIC;
                signal module_input33 :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal module_input42 :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal out_port_from_the_gpib_leds :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal out_port_from_the_gpio2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal out_port_from_the_led_pio :  STD_LOGIC;
                signal outputenable_n_to_the_ssram :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_debugaccess :  STD_LOGIC;
                signal pipeline_bridge_before_tristate_m1_endofpacket :  STD_LOGIC;
                signal pll_c2_out :  STD_LOGIC;
                signal pll_c3_out :  STD_LOGIC;
                signal read_n_to_the_cfi_flash :  STD_LOGIC;
                signal reset_n :  STD_LOGIC;
                signal reset_n_to_the_ssram :  STD_LOGIC;
                signal reset_phy_clk_n_from_the_ddr_sdram :  STD_LOGIC;
                signal select_n_to_the_cfi_flash :  STD_LOGIC;
                signal ssram_clk :  STD_LOGIC;
                signal write_n_to_the_cfi_flash :  STD_LOGIC;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your component and signal declaration here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


begin

  --Set us up the Dut
  DUT : gpib_edm1
    port map(
      MOSI_from_the_ad7928 => MOSI_from_the_ad7928,
      MOSI_from_the_dac_ad5308 => MOSI_from_the_dac_ad5308,
      SCLK_from_the_ad7928 => SCLK_from_the_ad7928,
      SCLK_from_the_dac_ad5308 => SCLK_from_the_dac_ad5308,
      SS_n_from_the_ad7928 => SS_n_from_the_ad7928,
      SS_n_from_the_dac_ad5308 => SS_n_from_the_dac_ad5308,
      adsc_n_to_the_ssram => adsc_n_to_the_ssram,
      bidir_port_to_and_from_the_gpio1 => bidir_port_to_and_from_the_gpio1,
      bw_n_to_the_ssram => bw_n_to_the_ssram,
      bwe_n_to_the_ssram => bwe_n_to_the_ssram,
      chipenable1_n_to_the_ssram => chipenable1_n_to_the_ssram,
      cpu_clk => cpu_clk,
      ddr_sdram_aux_full_rate_clk_out => ddr_sdram_aux_full_rate_clk_out,
      ddr_sdram_aux_half_rate_clk_out => ddr_sdram_aux_half_rate_clk_out,
      ddr_sdram_phy_clk_out => ddr_sdram_phy_clk_out,
      flash_ssram_tristate_address => flash_ssram_tristate_address,
      flash_ssram_tristate_data => flash_ssram_tristate_data,
      local_init_done_from_the_ddr_sdram => local_init_done_from_the_ddr_sdram,
      local_refresh_ack_from_the_ddr_sdram => local_refresh_ack_from_the_ddr_sdram,
      local_wdata_req_from_the_ddr_sdram => local_wdata_req_from_the_ddr_sdram,
      mem_addr_from_the_ddr_sdram => mem_addr_from_the_ddr_sdram,
      mem_ba_from_the_ddr_sdram => mem_ba_from_the_ddr_sdram,
      mem_cas_n_from_the_ddr_sdram => mem_cas_n_from_the_ddr_sdram,
      mem_cke_from_the_ddr_sdram => mem_cke_from_the_ddr_sdram,
      mem_clk_n_to_and_from_the_ddr_sdram => mem_clk_n_to_and_from_the_ddr_sdram,
      mem_clk_to_and_from_the_ddr_sdram => mem_clk_to_and_from_the_ddr_sdram,
      mem_cs_n_from_the_ddr_sdram => mem_cs_n_from_the_ddr_sdram,
      mem_dm_from_the_ddr_sdram => mem_dm_from_the_ddr_sdram,
      mem_dq_to_and_from_the_ddr_sdram => mem_dq_to_and_from_the_ddr_sdram,
      mem_dqs_to_and_from_the_ddr_sdram => mem_dqs_to_and_from_the_ddr_sdram,
      mem_ras_n_from_the_ddr_sdram => mem_ras_n_from_the_ddr_sdram,
      mem_we_n_from_the_ddr_sdram => mem_we_n_from_the_ddr_sdram,
      out_port_from_the_gpib_leds => out_port_from_the_gpib_leds,
      out_port_from_the_gpio2 => out_port_from_the_gpio2,
      out_port_from_the_led_pio => out_port_from_the_led_pio,
      outputenable_n_to_the_ssram => outputenable_n_to_the_ssram,
      pll_c2_out => pll_c2_out,
      pll_c3_out => pll_c3_out,
      read_n_to_the_cfi_flash => read_n_to_the_cfi_flash,
      reset_n_to_the_ssram => reset_n_to_the_ssram,
      reset_phy_clk_n_from_the_ddr_sdram => reset_phy_clk_n_from_the_ddr_sdram,
      select_n_to_the_cfi_flash => select_n_to_the_cfi_flash,
      ssram_clk => ssram_clk,
      write_n_to_the_cfi_flash => write_n_to_the_cfi_flash,
      MISO_to_the_ad7928 => MISO_to_the_ad7928,
      MISO_to_the_dac_ad5308 => MISO_to_the_dac_ad5308,
      clk_0 => clk_0,
      global_reset_n_to_the_ddr_sdram => global_reset_n_to_the_ddr_sdram,
      reset_n => reset_n
    );


  --the_cfi_flash, which is an e_ptf_instance
  the_cfi_flash : cfi_flash
    port map(
      data => flash_ssram_tristate_data (15 DOWNTO 0),
      address => module_input33,
      read_n => read_n_to_the_cfi_flash,
      select_n => select_n_to_the_cfi_flash,
      write_n => write_n_to_the_cfi_flash
    );

  module_input33 <= flash_ssram_tristate_address(23 DOWNTO 1);

  --the_ssram, which is an e_ptf_instance
  the_ssram : ssram
    port map(
      data => flash_ssram_tristate_data,
      address => module_input42,
      adsc_n => adsc_n_to_the_ssram,
      bw_n => bw_n_to_the_ssram,
      bwe_n => bwe_n_to_the_ssram,
      chipenable1_n => chipenable1_n_to_the_ssram,
      clk => cpu_clk,
      outputenable_n => outputenable_n_to_the_ssram,
      reset_n => reset_n_to_the_ssram
    );

  module_input42 <= flash_ssram_tristate_address(19 DOWNTO 2);

  process
  begin
    clk_0 <= '0';
    loop
       wait for 10 ns;
       clk_0 <= not clk_0;
    end loop;
  end process;
  PROCESS
    BEGIN
       reset_n <= '0';
       wait for 200 ns;
       reset_n <= '1'; 
    WAIT;
  END PROCESS;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add additional architecture here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


end europa;



--synthesis translate_on
